// Generator : SpinalHDL v1.12.3    git head : 591e64062329e5e2e2b81f4d52422948053edb97
// Component : SInt_ReuseC_SystolicArray_16x16
// Git hash  : 3085cb43943eb4f27ae7a21a20f2551c4c474ca1

`timescale 1ns/1ps

module SInt_ReuseC_SystolicArray_16x16 (
  input  wire [7:0]    io_inputA_0,
  input  wire [7:0]    io_inputA_1,
  input  wire [7:0]    io_inputA_2,
  input  wire [7:0]    io_inputA_3,
  input  wire [7:0]    io_inputA_4,
  input  wire [7:0]    io_inputA_5,
  input  wire [7:0]    io_inputA_6,
  input  wire [7:0]    io_inputA_7,
  input  wire [7:0]    io_inputA_8,
  input  wire [7:0]    io_inputA_9,
  input  wire [7:0]    io_inputA_10,
  input  wire [7:0]    io_inputA_11,
  input  wire [7:0]    io_inputA_12,
  input  wire [7:0]    io_inputA_13,
  input  wire [7:0]    io_inputA_14,
  input  wire [7:0]    io_inputA_15,
  input  wire [7:0]    io_inputB_0,
  input  wire [7:0]    io_inputB_1,
  input  wire [7:0]    io_inputB_2,
  input  wire [7:0]    io_inputB_3,
  input  wire [7:0]    io_inputB_4,
  input  wire [7:0]    io_inputB_5,
  input  wire [7:0]    io_inputB_6,
  input  wire [7:0]    io_inputB_7,
  input  wire [7:0]    io_inputB_8,
  input  wire [7:0]    io_inputB_9,
  input  wire [7:0]    io_inputB_10,
  input  wire [7:0]    io_inputB_11,
  input  wire [7:0]    io_inputB_12,
  input  wire [7:0]    io_inputB_13,
  input  wire [7:0]    io_inputB_14,
  input  wire [7:0]    io_inputB_15,
  input  wire          io_outputCaptureEnableC_0_0,
  input  wire          io_outputCaptureEnableC_0_1,
  input  wire          io_outputCaptureEnableC_0_2,
  input  wire          io_outputCaptureEnableC_0_3,
  input  wire          io_outputCaptureEnableC_0_4,
  input  wire          io_outputCaptureEnableC_0_5,
  input  wire          io_outputCaptureEnableC_0_6,
  input  wire          io_outputCaptureEnableC_0_7,
  input  wire          io_outputCaptureEnableC_0_8,
  input  wire          io_outputCaptureEnableC_0_9,
  input  wire          io_outputCaptureEnableC_0_10,
  input  wire          io_outputCaptureEnableC_0_11,
  input  wire          io_outputCaptureEnableC_0_12,
  input  wire          io_outputCaptureEnableC_0_13,
  input  wire          io_outputCaptureEnableC_0_14,
  input  wire          io_outputCaptureEnableC_0_15,
  input  wire          io_outputCaptureEnableC_1_0,
  input  wire          io_outputCaptureEnableC_1_1,
  input  wire          io_outputCaptureEnableC_1_2,
  input  wire          io_outputCaptureEnableC_1_3,
  input  wire          io_outputCaptureEnableC_1_4,
  input  wire          io_outputCaptureEnableC_1_5,
  input  wire          io_outputCaptureEnableC_1_6,
  input  wire          io_outputCaptureEnableC_1_7,
  input  wire          io_outputCaptureEnableC_1_8,
  input  wire          io_outputCaptureEnableC_1_9,
  input  wire          io_outputCaptureEnableC_1_10,
  input  wire          io_outputCaptureEnableC_1_11,
  input  wire          io_outputCaptureEnableC_1_12,
  input  wire          io_outputCaptureEnableC_1_13,
  input  wire          io_outputCaptureEnableC_1_14,
  input  wire          io_outputCaptureEnableC_1_15,
  input  wire          io_outputCaptureEnableC_2_0,
  input  wire          io_outputCaptureEnableC_2_1,
  input  wire          io_outputCaptureEnableC_2_2,
  input  wire          io_outputCaptureEnableC_2_3,
  input  wire          io_outputCaptureEnableC_2_4,
  input  wire          io_outputCaptureEnableC_2_5,
  input  wire          io_outputCaptureEnableC_2_6,
  input  wire          io_outputCaptureEnableC_2_7,
  input  wire          io_outputCaptureEnableC_2_8,
  input  wire          io_outputCaptureEnableC_2_9,
  input  wire          io_outputCaptureEnableC_2_10,
  input  wire          io_outputCaptureEnableC_2_11,
  input  wire          io_outputCaptureEnableC_2_12,
  input  wire          io_outputCaptureEnableC_2_13,
  input  wire          io_outputCaptureEnableC_2_14,
  input  wire          io_outputCaptureEnableC_2_15,
  input  wire          io_outputCaptureEnableC_3_0,
  input  wire          io_outputCaptureEnableC_3_1,
  input  wire          io_outputCaptureEnableC_3_2,
  input  wire          io_outputCaptureEnableC_3_3,
  input  wire          io_outputCaptureEnableC_3_4,
  input  wire          io_outputCaptureEnableC_3_5,
  input  wire          io_outputCaptureEnableC_3_6,
  input  wire          io_outputCaptureEnableC_3_7,
  input  wire          io_outputCaptureEnableC_3_8,
  input  wire          io_outputCaptureEnableC_3_9,
  input  wire          io_outputCaptureEnableC_3_10,
  input  wire          io_outputCaptureEnableC_3_11,
  input  wire          io_outputCaptureEnableC_3_12,
  input  wire          io_outputCaptureEnableC_3_13,
  input  wire          io_outputCaptureEnableC_3_14,
  input  wire          io_outputCaptureEnableC_3_15,
  input  wire          io_outputCaptureEnableC_4_0,
  input  wire          io_outputCaptureEnableC_4_1,
  input  wire          io_outputCaptureEnableC_4_2,
  input  wire          io_outputCaptureEnableC_4_3,
  input  wire          io_outputCaptureEnableC_4_4,
  input  wire          io_outputCaptureEnableC_4_5,
  input  wire          io_outputCaptureEnableC_4_6,
  input  wire          io_outputCaptureEnableC_4_7,
  input  wire          io_outputCaptureEnableC_4_8,
  input  wire          io_outputCaptureEnableC_4_9,
  input  wire          io_outputCaptureEnableC_4_10,
  input  wire          io_outputCaptureEnableC_4_11,
  input  wire          io_outputCaptureEnableC_4_12,
  input  wire          io_outputCaptureEnableC_4_13,
  input  wire          io_outputCaptureEnableC_4_14,
  input  wire          io_outputCaptureEnableC_4_15,
  input  wire          io_outputCaptureEnableC_5_0,
  input  wire          io_outputCaptureEnableC_5_1,
  input  wire          io_outputCaptureEnableC_5_2,
  input  wire          io_outputCaptureEnableC_5_3,
  input  wire          io_outputCaptureEnableC_5_4,
  input  wire          io_outputCaptureEnableC_5_5,
  input  wire          io_outputCaptureEnableC_5_6,
  input  wire          io_outputCaptureEnableC_5_7,
  input  wire          io_outputCaptureEnableC_5_8,
  input  wire          io_outputCaptureEnableC_5_9,
  input  wire          io_outputCaptureEnableC_5_10,
  input  wire          io_outputCaptureEnableC_5_11,
  input  wire          io_outputCaptureEnableC_5_12,
  input  wire          io_outputCaptureEnableC_5_13,
  input  wire          io_outputCaptureEnableC_5_14,
  input  wire          io_outputCaptureEnableC_5_15,
  input  wire          io_outputCaptureEnableC_6_0,
  input  wire          io_outputCaptureEnableC_6_1,
  input  wire          io_outputCaptureEnableC_6_2,
  input  wire          io_outputCaptureEnableC_6_3,
  input  wire          io_outputCaptureEnableC_6_4,
  input  wire          io_outputCaptureEnableC_6_5,
  input  wire          io_outputCaptureEnableC_6_6,
  input  wire          io_outputCaptureEnableC_6_7,
  input  wire          io_outputCaptureEnableC_6_8,
  input  wire          io_outputCaptureEnableC_6_9,
  input  wire          io_outputCaptureEnableC_6_10,
  input  wire          io_outputCaptureEnableC_6_11,
  input  wire          io_outputCaptureEnableC_6_12,
  input  wire          io_outputCaptureEnableC_6_13,
  input  wire          io_outputCaptureEnableC_6_14,
  input  wire          io_outputCaptureEnableC_6_15,
  input  wire          io_outputCaptureEnableC_7_0,
  input  wire          io_outputCaptureEnableC_7_1,
  input  wire          io_outputCaptureEnableC_7_2,
  input  wire          io_outputCaptureEnableC_7_3,
  input  wire          io_outputCaptureEnableC_7_4,
  input  wire          io_outputCaptureEnableC_7_5,
  input  wire          io_outputCaptureEnableC_7_6,
  input  wire          io_outputCaptureEnableC_7_7,
  input  wire          io_outputCaptureEnableC_7_8,
  input  wire          io_outputCaptureEnableC_7_9,
  input  wire          io_outputCaptureEnableC_7_10,
  input  wire          io_outputCaptureEnableC_7_11,
  input  wire          io_outputCaptureEnableC_7_12,
  input  wire          io_outputCaptureEnableC_7_13,
  input  wire          io_outputCaptureEnableC_7_14,
  input  wire          io_outputCaptureEnableC_7_15,
  input  wire          io_outputCaptureEnableC_8_0,
  input  wire          io_outputCaptureEnableC_8_1,
  input  wire          io_outputCaptureEnableC_8_2,
  input  wire          io_outputCaptureEnableC_8_3,
  input  wire          io_outputCaptureEnableC_8_4,
  input  wire          io_outputCaptureEnableC_8_5,
  input  wire          io_outputCaptureEnableC_8_6,
  input  wire          io_outputCaptureEnableC_8_7,
  input  wire          io_outputCaptureEnableC_8_8,
  input  wire          io_outputCaptureEnableC_8_9,
  input  wire          io_outputCaptureEnableC_8_10,
  input  wire          io_outputCaptureEnableC_8_11,
  input  wire          io_outputCaptureEnableC_8_12,
  input  wire          io_outputCaptureEnableC_8_13,
  input  wire          io_outputCaptureEnableC_8_14,
  input  wire          io_outputCaptureEnableC_8_15,
  input  wire          io_outputCaptureEnableC_9_0,
  input  wire          io_outputCaptureEnableC_9_1,
  input  wire          io_outputCaptureEnableC_9_2,
  input  wire          io_outputCaptureEnableC_9_3,
  input  wire          io_outputCaptureEnableC_9_4,
  input  wire          io_outputCaptureEnableC_9_5,
  input  wire          io_outputCaptureEnableC_9_6,
  input  wire          io_outputCaptureEnableC_9_7,
  input  wire          io_outputCaptureEnableC_9_8,
  input  wire          io_outputCaptureEnableC_9_9,
  input  wire          io_outputCaptureEnableC_9_10,
  input  wire          io_outputCaptureEnableC_9_11,
  input  wire          io_outputCaptureEnableC_9_12,
  input  wire          io_outputCaptureEnableC_9_13,
  input  wire          io_outputCaptureEnableC_9_14,
  input  wire          io_outputCaptureEnableC_9_15,
  input  wire          io_outputCaptureEnableC_10_0,
  input  wire          io_outputCaptureEnableC_10_1,
  input  wire          io_outputCaptureEnableC_10_2,
  input  wire          io_outputCaptureEnableC_10_3,
  input  wire          io_outputCaptureEnableC_10_4,
  input  wire          io_outputCaptureEnableC_10_5,
  input  wire          io_outputCaptureEnableC_10_6,
  input  wire          io_outputCaptureEnableC_10_7,
  input  wire          io_outputCaptureEnableC_10_8,
  input  wire          io_outputCaptureEnableC_10_9,
  input  wire          io_outputCaptureEnableC_10_10,
  input  wire          io_outputCaptureEnableC_10_11,
  input  wire          io_outputCaptureEnableC_10_12,
  input  wire          io_outputCaptureEnableC_10_13,
  input  wire          io_outputCaptureEnableC_10_14,
  input  wire          io_outputCaptureEnableC_10_15,
  input  wire          io_outputCaptureEnableC_11_0,
  input  wire          io_outputCaptureEnableC_11_1,
  input  wire          io_outputCaptureEnableC_11_2,
  input  wire          io_outputCaptureEnableC_11_3,
  input  wire          io_outputCaptureEnableC_11_4,
  input  wire          io_outputCaptureEnableC_11_5,
  input  wire          io_outputCaptureEnableC_11_6,
  input  wire          io_outputCaptureEnableC_11_7,
  input  wire          io_outputCaptureEnableC_11_8,
  input  wire          io_outputCaptureEnableC_11_9,
  input  wire          io_outputCaptureEnableC_11_10,
  input  wire          io_outputCaptureEnableC_11_11,
  input  wire          io_outputCaptureEnableC_11_12,
  input  wire          io_outputCaptureEnableC_11_13,
  input  wire          io_outputCaptureEnableC_11_14,
  input  wire          io_outputCaptureEnableC_11_15,
  input  wire          io_outputCaptureEnableC_12_0,
  input  wire          io_outputCaptureEnableC_12_1,
  input  wire          io_outputCaptureEnableC_12_2,
  input  wire          io_outputCaptureEnableC_12_3,
  input  wire          io_outputCaptureEnableC_12_4,
  input  wire          io_outputCaptureEnableC_12_5,
  input  wire          io_outputCaptureEnableC_12_6,
  input  wire          io_outputCaptureEnableC_12_7,
  input  wire          io_outputCaptureEnableC_12_8,
  input  wire          io_outputCaptureEnableC_12_9,
  input  wire          io_outputCaptureEnableC_12_10,
  input  wire          io_outputCaptureEnableC_12_11,
  input  wire          io_outputCaptureEnableC_12_12,
  input  wire          io_outputCaptureEnableC_12_13,
  input  wire          io_outputCaptureEnableC_12_14,
  input  wire          io_outputCaptureEnableC_12_15,
  input  wire          io_outputCaptureEnableC_13_0,
  input  wire          io_outputCaptureEnableC_13_1,
  input  wire          io_outputCaptureEnableC_13_2,
  input  wire          io_outputCaptureEnableC_13_3,
  input  wire          io_outputCaptureEnableC_13_4,
  input  wire          io_outputCaptureEnableC_13_5,
  input  wire          io_outputCaptureEnableC_13_6,
  input  wire          io_outputCaptureEnableC_13_7,
  input  wire          io_outputCaptureEnableC_13_8,
  input  wire          io_outputCaptureEnableC_13_9,
  input  wire          io_outputCaptureEnableC_13_10,
  input  wire          io_outputCaptureEnableC_13_11,
  input  wire          io_outputCaptureEnableC_13_12,
  input  wire          io_outputCaptureEnableC_13_13,
  input  wire          io_outputCaptureEnableC_13_14,
  input  wire          io_outputCaptureEnableC_13_15,
  input  wire          io_outputCaptureEnableC_14_0,
  input  wire          io_outputCaptureEnableC_14_1,
  input  wire          io_outputCaptureEnableC_14_2,
  input  wire          io_outputCaptureEnableC_14_3,
  input  wire          io_outputCaptureEnableC_14_4,
  input  wire          io_outputCaptureEnableC_14_5,
  input  wire          io_outputCaptureEnableC_14_6,
  input  wire          io_outputCaptureEnableC_14_7,
  input  wire          io_outputCaptureEnableC_14_8,
  input  wire          io_outputCaptureEnableC_14_9,
  input  wire          io_outputCaptureEnableC_14_10,
  input  wire          io_outputCaptureEnableC_14_11,
  input  wire          io_outputCaptureEnableC_14_12,
  input  wire          io_outputCaptureEnableC_14_13,
  input  wire          io_outputCaptureEnableC_14_14,
  input  wire          io_outputCaptureEnableC_14_15,
  input  wire          io_outputCaptureEnableC_15_0,
  input  wire          io_outputCaptureEnableC_15_1,
  input  wire          io_outputCaptureEnableC_15_2,
  input  wire          io_outputCaptureEnableC_15_3,
  input  wire          io_outputCaptureEnableC_15_4,
  input  wire          io_outputCaptureEnableC_15_5,
  input  wire          io_outputCaptureEnableC_15_6,
  input  wire          io_outputCaptureEnableC_15_7,
  input  wire          io_outputCaptureEnableC_15_8,
  input  wire          io_outputCaptureEnableC_15_9,
  input  wire          io_outputCaptureEnableC_15_10,
  input  wire          io_outputCaptureEnableC_15_11,
  input  wire          io_outputCaptureEnableC_15_12,
  input  wire          io_outputCaptureEnableC_15_13,
  input  wire          io_outputCaptureEnableC_15_14,
  input  wire          io_outputCaptureEnableC_15_15,
  input  wire          io_resetPartialC_0_0,
  input  wire          io_resetPartialC_0_1,
  input  wire          io_resetPartialC_0_2,
  input  wire          io_resetPartialC_0_3,
  input  wire          io_resetPartialC_0_4,
  input  wire          io_resetPartialC_0_5,
  input  wire          io_resetPartialC_0_6,
  input  wire          io_resetPartialC_0_7,
  input  wire          io_resetPartialC_0_8,
  input  wire          io_resetPartialC_0_9,
  input  wire          io_resetPartialC_0_10,
  input  wire          io_resetPartialC_0_11,
  input  wire          io_resetPartialC_0_12,
  input  wire          io_resetPartialC_0_13,
  input  wire          io_resetPartialC_0_14,
  input  wire          io_resetPartialC_0_15,
  input  wire          io_resetPartialC_1_0,
  input  wire          io_resetPartialC_1_1,
  input  wire          io_resetPartialC_1_2,
  input  wire          io_resetPartialC_1_3,
  input  wire          io_resetPartialC_1_4,
  input  wire          io_resetPartialC_1_5,
  input  wire          io_resetPartialC_1_6,
  input  wire          io_resetPartialC_1_7,
  input  wire          io_resetPartialC_1_8,
  input  wire          io_resetPartialC_1_9,
  input  wire          io_resetPartialC_1_10,
  input  wire          io_resetPartialC_1_11,
  input  wire          io_resetPartialC_1_12,
  input  wire          io_resetPartialC_1_13,
  input  wire          io_resetPartialC_1_14,
  input  wire          io_resetPartialC_1_15,
  input  wire          io_resetPartialC_2_0,
  input  wire          io_resetPartialC_2_1,
  input  wire          io_resetPartialC_2_2,
  input  wire          io_resetPartialC_2_3,
  input  wire          io_resetPartialC_2_4,
  input  wire          io_resetPartialC_2_5,
  input  wire          io_resetPartialC_2_6,
  input  wire          io_resetPartialC_2_7,
  input  wire          io_resetPartialC_2_8,
  input  wire          io_resetPartialC_2_9,
  input  wire          io_resetPartialC_2_10,
  input  wire          io_resetPartialC_2_11,
  input  wire          io_resetPartialC_2_12,
  input  wire          io_resetPartialC_2_13,
  input  wire          io_resetPartialC_2_14,
  input  wire          io_resetPartialC_2_15,
  input  wire          io_resetPartialC_3_0,
  input  wire          io_resetPartialC_3_1,
  input  wire          io_resetPartialC_3_2,
  input  wire          io_resetPartialC_3_3,
  input  wire          io_resetPartialC_3_4,
  input  wire          io_resetPartialC_3_5,
  input  wire          io_resetPartialC_3_6,
  input  wire          io_resetPartialC_3_7,
  input  wire          io_resetPartialC_3_8,
  input  wire          io_resetPartialC_3_9,
  input  wire          io_resetPartialC_3_10,
  input  wire          io_resetPartialC_3_11,
  input  wire          io_resetPartialC_3_12,
  input  wire          io_resetPartialC_3_13,
  input  wire          io_resetPartialC_3_14,
  input  wire          io_resetPartialC_3_15,
  input  wire          io_resetPartialC_4_0,
  input  wire          io_resetPartialC_4_1,
  input  wire          io_resetPartialC_4_2,
  input  wire          io_resetPartialC_4_3,
  input  wire          io_resetPartialC_4_4,
  input  wire          io_resetPartialC_4_5,
  input  wire          io_resetPartialC_4_6,
  input  wire          io_resetPartialC_4_7,
  input  wire          io_resetPartialC_4_8,
  input  wire          io_resetPartialC_4_9,
  input  wire          io_resetPartialC_4_10,
  input  wire          io_resetPartialC_4_11,
  input  wire          io_resetPartialC_4_12,
  input  wire          io_resetPartialC_4_13,
  input  wire          io_resetPartialC_4_14,
  input  wire          io_resetPartialC_4_15,
  input  wire          io_resetPartialC_5_0,
  input  wire          io_resetPartialC_5_1,
  input  wire          io_resetPartialC_5_2,
  input  wire          io_resetPartialC_5_3,
  input  wire          io_resetPartialC_5_4,
  input  wire          io_resetPartialC_5_5,
  input  wire          io_resetPartialC_5_6,
  input  wire          io_resetPartialC_5_7,
  input  wire          io_resetPartialC_5_8,
  input  wire          io_resetPartialC_5_9,
  input  wire          io_resetPartialC_5_10,
  input  wire          io_resetPartialC_5_11,
  input  wire          io_resetPartialC_5_12,
  input  wire          io_resetPartialC_5_13,
  input  wire          io_resetPartialC_5_14,
  input  wire          io_resetPartialC_5_15,
  input  wire          io_resetPartialC_6_0,
  input  wire          io_resetPartialC_6_1,
  input  wire          io_resetPartialC_6_2,
  input  wire          io_resetPartialC_6_3,
  input  wire          io_resetPartialC_6_4,
  input  wire          io_resetPartialC_6_5,
  input  wire          io_resetPartialC_6_6,
  input  wire          io_resetPartialC_6_7,
  input  wire          io_resetPartialC_6_8,
  input  wire          io_resetPartialC_6_9,
  input  wire          io_resetPartialC_6_10,
  input  wire          io_resetPartialC_6_11,
  input  wire          io_resetPartialC_6_12,
  input  wire          io_resetPartialC_6_13,
  input  wire          io_resetPartialC_6_14,
  input  wire          io_resetPartialC_6_15,
  input  wire          io_resetPartialC_7_0,
  input  wire          io_resetPartialC_7_1,
  input  wire          io_resetPartialC_7_2,
  input  wire          io_resetPartialC_7_3,
  input  wire          io_resetPartialC_7_4,
  input  wire          io_resetPartialC_7_5,
  input  wire          io_resetPartialC_7_6,
  input  wire          io_resetPartialC_7_7,
  input  wire          io_resetPartialC_7_8,
  input  wire          io_resetPartialC_7_9,
  input  wire          io_resetPartialC_7_10,
  input  wire          io_resetPartialC_7_11,
  input  wire          io_resetPartialC_7_12,
  input  wire          io_resetPartialC_7_13,
  input  wire          io_resetPartialC_7_14,
  input  wire          io_resetPartialC_7_15,
  input  wire          io_resetPartialC_8_0,
  input  wire          io_resetPartialC_8_1,
  input  wire          io_resetPartialC_8_2,
  input  wire          io_resetPartialC_8_3,
  input  wire          io_resetPartialC_8_4,
  input  wire          io_resetPartialC_8_5,
  input  wire          io_resetPartialC_8_6,
  input  wire          io_resetPartialC_8_7,
  input  wire          io_resetPartialC_8_8,
  input  wire          io_resetPartialC_8_9,
  input  wire          io_resetPartialC_8_10,
  input  wire          io_resetPartialC_8_11,
  input  wire          io_resetPartialC_8_12,
  input  wire          io_resetPartialC_8_13,
  input  wire          io_resetPartialC_8_14,
  input  wire          io_resetPartialC_8_15,
  input  wire          io_resetPartialC_9_0,
  input  wire          io_resetPartialC_9_1,
  input  wire          io_resetPartialC_9_2,
  input  wire          io_resetPartialC_9_3,
  input  wire          io_resetPartialC_9_4,
  input  wire          io_resetPartialC_9_5,
  input  wire          io_resetPartialC_9_6,
  input  wire          io_resetPartialC_9_7,
  input  wire          io_resetPartialC_9_8,
  input  wire          io_resetPartialC_9_9,
  input  wire          io_resetPartialC_9_10,
  input  wire          io_resetPartialC_9_11,
  input  wire          io_resetPartialC_9_12,
  input  wire          io_resetPartialC_9_13,
  input  wire          io_resetPartialC_9_14,
  input  wire          io_resetPartialC_9_15,
  input  wire          io_resetPartialC_10_0,
  input  wire          io_resetPartialC_10_1,
  input  wire          io_resetPartialC_10_2,
  input  wire          io_resetPartialC_10_3,
  input  wire          io_resetPartialC_10_4,
  input  wire          io_resetPartialC_10_5,
  input  wire          io_resetPartialC_10_6,
  input  wire          io_resetPartialC_10_7,
  input  wire          io_resetPartialC_10_8,
  input  wire          io_resetPartialC_10_9,
  input  wire          io_resetPartialC_10_10,
  input  wire          io_resetPartialC_10_11,
  input  wire          io_resetPartialC_10_12,
  input  wire          io_resetPartialC_10_13,
  input  wire          io_resetPartialC_10_14,
  input  wire          io_resetPartialC_10_15,
  input  wire          io_resetPartialC_11_0,
  input  wire          io_resetPartialC_11_1,
  input  wire          io_resetPartialC_11_2,
  input  wire          io_resetPartialC_11_3,
  input  wire          io_resetPartialC_11_4,
  input  wire          io_resetPartialC_11_5,
  input  wire          io_resetPartialC_11_6,
  input  wire          io_resetPartialC_11_7,
  input  wire          io_resetPartialC_11_8,
  input  wire          io_resetPartialC_11_9,
  input  wire          io_resetPartialC_11_10,
  input  wire          io_resetPartialC_11_11,
  input  wire          io_resetPartialC_11_12,
  input  wire          io_resetPartialC_11_13,
  input  wire          io_resetPartialC_11_14,
  input  wire          io_resetPartialC_11_15,
  input  wire          io_resetPartialC_12_0,
  input  wire          io_resetPartialC_12_1,
  input  wire          io_resetPartialC_12_2,
  input  wire          io_resetPartialC_12_3,
  input  wire          io_resetPartialC_12_4,
  input  wire          io_resetPartialC_12_5,
  input  wire          io_resetPartialC_12_6,
  input  wire          io_resetPartialC_12_7,
  input  wire          io_resetPartialC_12_8,
  input  wire          io_resetPartialC_12_9,
  input  wire          io_resetPartialC_12_10,
  input  wire          io_resetPartialC_12_11,
  input  wire          io_resetPartialC_12_12,
  input  wire          io_resetPartialC_12_13,
  input  wire          io_resetPartialC_12_14,
  input  wire          io_resetPartialC_12_15,
  input  wire          io_resetPartialC_13_0,
  input  wire          io_resetPartialC_13_1,
  input  wire          io_resetPartialC_13_2,
  input  wire          io_resetPartialC_13_3,
  input  wire          io_resetPartialC_13_4,
  input  wire          io_resetPartialC_13_5,
  input  wire          io_resetPartialC_13_6,
  input  wire          io_resetPartialC_13_7,
  input  wire          io_resetPartialC_13_8,
  input  wire          io_resetPartialC_13_9,
  input  wire          io_resetPartialC_13_10,
  input  wire          io_resetPartialC_13_11,
  input  wire          io_resetPartialC_13_12,
  input  wire          io_resetPartialC_13_13,
  input  wire          io_resetPartialC_13_14,
  input  wire          io_resetPartialC_13_15,
  input  wire          io_resetPartialC_14_0,
  input  wire          io_resetPartialC_14_1,
  input  wire          io_resetPartialC_14_2,
  input  wire          io_resetPartialC_14_3,
  input  wire          io_resetPartialC_14_4,
  input  wire          io_resetPartialC_14_5,
  input  wire          io_resetPartialC_14_6,
  input  wire          io_resetPartialC_14_7,
  input  wire          io_resetPartialC_14_8,
  input  wire          io_resetPartialC_14_9,
  input  wire          io_resetPartialC_14_10,
  input  wire          io_resetPartialC_14_11,
  input  wire          io_resetPartialC_14_12,
  input  wire          io_resetPartialC_14_13,
  input  wire          io_resetPartialC_14_14,
  input  wire          io_resetPartialC_14_15,
  input  wire          io_resetPartialC_15_0,
  input  wire          io_resetPartialC_15_1,
  input  wire          io_resetPartialC_15_2,
  input  wire          io_resetPartialC_15_3,
  input  wire          io_resetPartialC_15_4,
  input  wire          io_resetPartialC_15_5,
  input  wire          io_resetPartialC_15_6,
  input  wire          io_resetPartialC_15_7,
  input  wire          io_resetPartialC_15_8,
  input  wire          io_resetPartialC_15_9,
  input  wire          io_resetPartialC_15_10,
  input  wire          io_resetPartialC_15_11,
  input  wire          io_resetPartialC_15_12,
  input  wire          io_resetPartialC_15_13,
  input  wire          io_resetPartialC_15_14,
  input  wire          io_resetPartialC_15_15,
  output wire [25:0]   io_outputC_0,
  output wire [25:0]   io_outputC_1,
  output wire [25:0]   io_outputC_2,
  output wire [25:0]   io_outputC_3,
  output wire [25:0]   io_outputC_4,
  output wire [25:0]   io_outputC_5,
  output wire [25:0]   io_outputC_6,
  output wire [25:0]   io_outputC_7,
  output wire [25:0]   io_outputC_8,
  output wire [25:0]   io_outputC_9,
  output wire [25:0]   io_outputC_10,
  output wire [25:0]   io_outputC_11,
  output wire [25:0]   io_outputC_12,
  output wire [25:0]   io_outputC_13,
  output wire [25:0]   io_outputC_14,
  output wire [25:0]   io_outputC_15,
  output wire [25:0]   io_outputC_16,
  output wire [25:0]   io_outputC_17,
  output wire [25:0]   io_outputC_18,
  output wire [25:0]   io_outputC_19,
  output wire [25:0]   io_outputC_20,
  output wire [25:0]   io_outputC_21,
  output wire [25:0]   io_outputC_22,
  output wire [25:0]   io_outputC_23,
  output wire [25:0]   io_outputC_24,
  output wire [25:0]   io_outputC_25,
  output wire [25:0]   io_outputC_26,
  output wire [25:0]   io_outputC_27,
  output wire [25:0]   io_outputC_28,
  output wire [25:0]   io_outputC_29,
  output wire [25:0]   io_outputC_30,
  input  wire          clk,
  input  wire          reset
);

  wire       [7:0]    pes_0_0_io_outputA;
  wire       [7:0]    pes_0_0_io_outputB;
  wire       [25:0]   pes_0_0_io_outputC;
  wire       [7:0]    pes_0_1_io_outputA;
  wire       [7:0]    pes_0_1_io_outputB;
  wire       [25:0]   pes_0_1_io_outputC;
  wire       [7:0]    pes_0_2_io_outputA;
  wire       [7:0]    pes_0_2_io_outputB;
  wire       [25:0]   pes_0_2_io_outputC;
  wire       [7:0]    pes_0_3_io_outputA;
  wire       [7:0]    pes_0_3_io_outputB;
  wire       [25:0]   pes_0_3_io_outputC;
  wire       [7:0]    pes_0_4_io_outputA;
  wire       [7:0]    pes_0_4_io_outputB;
  wire       [25:0]   pes_0_4_io_outputC;
  wire       [7:0]    pes_0_5_io_outputA;
  wire       [7:0]    pes_0_5_io_outputB;
  wire       [25:0]   pes_0_5_io_outputC;
  wire       [7:0]    pes_0_6_io_outputA;
  wire       [7:0]    pes_0_6_io_outputB;
  wire       [25:0]   pes_0_6_io_outputC;
  wire       [7:0]    pes_0_7_io_outputA;
  wire       [7:0]    pes_0_7_io_outputB;
  wire       [25:0]   pes_0_7_io_outputC;
  wire       [7:0]    pes_0_8_io_outputA;
  wire       [7:0]    pes_0_8_io_outputB;
  wire       [25:0]   pes_0_8_io_outputC;
  wire       [7:0]    pes_0_9_io_outputA;
  wire       [7:0]    pes_0_9_io_outputB;
  wire       [25:0]   pes_0_9_io_outputC;
  wire       [7:0]    pes_0_10_io_outputA;
  wire       [7:0]    pes_0_10_io_outputB;
  wire       [25:0]   pes_0_10_io_outputC;
  wire       [7:0]    pes_0_11_io_outputA;
  wire       [7:0]    pes_0_11_io_outputB;
  wire       [25:0]   pes_0_11_io_outputC;
  wire       [7:0]    pes_0_12_io_outputA;
  wire       [7:0]    pes_0_12_io_outputB;
  wire       [25:0]   pes_0_12_io_outputC;
  wire       [7:0]    pes_0_13_io_outputA;
  wire       [7:0]    pes_0_13_io_outputB;
  wire       [25:0]   pes_0_13_io_outputC;
  wire       [7:0]    pes_0_14_io_outputA;
  wire       [7:0]    pes_0_14_io_outputB;
  wire       [25:0]   pes_0_14_io_outputC;
  wire       [7:0]    pes_0_15_io_outputB;
  wire       [25:0]   pes_0_15_io_outputC;
  wire       [7:0]    pes_1_0_io_outputA;
  wire       [7:0]    pes_1_0_io_outputB;
  wire       [25:0]   pes_1_0_io_outputC;
  wire       [7:0]    pes_1_1_io_outputA;
  wire       [7:0]    pes_1_1_io_outputB;
  wire       [25:0]   pes_1_1_io_outputC;
  wire       [7:0]    pes_1_2_io_outputA;
  wire       [7:0]    pes_1_2_io_outputB;
  wire       [25:0]   pes_1_2_io_outputC;
  wire       [7:0]    pes_1_3_io_outputA;
  wire       [7:0]    pes_1_3_io_outputB;
  wire       [25:0]   pes_1_3_io_outputC;
  wire       [7:0]    pes_1_4_io_outputA;
  wire       [7:0]    pes_1_4_io_outputB;
  wire       [25:0]   pes_1_4_io_outputC;
  wire       [7:0]    pes_1_5_io_outputA;
  wire       [7:0]    pes_1_5_io_outputB;
  wire       [25:0]   pes_1_5_io_outputC;
  wire       [7:0]    pes_1_6_io_outputA;
  wire       [7:0]    pes_1_6_io_outputB;
  wire       [25:0]   pes_1_6_io_outputC;
  wire       [7:0]    pes_1_7_io_outputA;
  wire       [7:0]    pes_1_7_io_outputB;
  wire       [25:0]   pes_1_7_io_outputC;
  wire       [7:0]    pes_1_8_io_outputA;
  wire       [7:0]    pes_1_8_io_outputB;
  wire       [25:0]   pes_1_8_io_outputC;
  wire       [7:0]    pes_1_9_io_outputA;
  wire       [7:0]    pes_1_9_io_outputB;
  wire       [25:0]   pes_1_9_io_outputC;
  wire       [7:0]    pes_1_10_io_outputA;
  wire       [7:0]    pes_1_10_io_outputB;
  wire       [25:0]   pes_1_10_io_outputC;
  wire       [7:0]    pes_1_11_io_outputA;
  wire       [7:0]    pes_1_11_io_outputB;
  wire       [25:0]   pes_1_11_io_outputC;
  wire       [7:0]    pes_1_12_io_outputA;
  wire       [7:0]    pes_1_12_io_outputB;
  wire       [25:0]   pes_1_12_io_outputC;
  wire       [7:0]    pes_1_13_io_outputA;
  wire       [7:0]    pes_1_13_io_outputB;
  wire       [25:0]   pes_1_13_io_outputC;
  wire       [7:0]    pes_1_14_io_outputA;
  wire       [7:0]    pes_1_14_io_outputB;
  wire       [25:0]   pes_1_14_io_outputC;
  wire       [7:0]    pes_1_15_io_outputB;
  wire       [25:0]   pes_1_15_io_outputC;
  wire       [7:0]    pes_2_0_io_outputA;
  wire       [7:0]    pes_2_0_io_outputB;
  wire       [25:0]   pes_2_0_io_outputC;
  wire       [7:0]    pes_2_1_io_outputA;
  wire       [7:0]    pes_2_1_io_outputB;
  wire       [25:0]   pes_2_1_io_outputC;
  wire       [7:0]    pes_2_2_io_outputA;
  wire       [7:0]    pes_2_2_io_outputB;
  wire       [25:0]   pes_2_2_io_outputC;
  wire       [7:0]    pes_2_3_io_outputA;
  wire       [7:0]    pes_2_3_io_outputB;
  wire       [25:0]   pes_2_3_io_outputC;
  wire       [7:0]    pes_2_4_io_outputA;
  wire       [7:0]    pes_2_4_io_outputB;
  wire       [25:0]   pes_2_4_io_outputC;
  wire       [7:0]    pes_2_5_io_outputA;
  wire       [7:0]    pes_2_5_io_outputB;
  wire       [25:0]   pes_2_5_io_outputC;
  wire       [7:0]    pes_2_6_io_outputA;
  wire       [7:0]    pes_2_6_io_outputB;
  wire       [25:0]   pes_2_6_io_outputC;
  wire       [7:0]    pes_2_7_io_outputA;
  wire       [7:0]    pes_2_7_io_outputB;
  wire       [25:0]   pes_2_7_io_outputC;
  wire       [7:0]    pes_2_8_io_outputA;
  wire       [7:0]    pes_2_8_io_outputB;
  wire       [25:0]   pes_2_8_io_outputC;
  wire       [7:0]    pes_2_9_io_outputA;
  wire       [7:0]    pes_2_9_io_outputB;
  wire       [25:0]   pes_2_9_io_outputC;
  wire       [7:0]    pes_2_10_io_outputA;
  wire       [7:0]    pes_2_10_io_outputB;
  wire       [25:0]   pes_2_10_io_outputC;
  wire       [7:0]    pes_2_11_io_outputA;
  wire       [7:0]    pes_2_11_io_outputB;
  wire       [25:0]   pes_2_11_io_outputC;
  wire       [7:0]    pes_2_12_io_outputA;
  wire       [7:0]    pes_2_12_io_outputB;
  wire       [25:0]   pes_2_12_io_outputC;
  wire       [7:0]    pes_2_13_io_outputA;
  wire       [7:0]    pes_2_13_io_outputB;
  wire       [25:0]   pes_2_13_io_outputC;
  wire       [7:0]    pes_2_14_io_outputA;
  wire       [7:0]    pes_2_14_io_outputB;
  wire       [25:0]   pes_2_14_io_outputC;
  wire       [7:0]    pes_2_15_io_outputB;
  wire       [25:0]   pes_2_15_io_outputC;
  wire       [7:0]    pes_3_0_io_outputA;
  wire       [7:0]    pes_3_0_io_outputB;
  wire       [25:0]   pes_3_0_io_outputC;
  wire       [7:0]    pes_3_1_io_outputA;
  wire       [7:0]    pes_3_1_io_outputB;
  wire       [25:0]   pes_3_1_io_outputC;
  wire       [7:0]    pes_3_2_io_outputA;
  wire       [7:0]    pes_3_2_io_outputB;
  wire       [25:0]   pes_3_2_io_outputC;
  wire       [7:0]    pes_3_3_io_outputA;
  wire       [7:0]    pes_3_3_io_outputB;
  wire       [25:0]   pes_3_3_io_outputC;
  wire       [7:0]    pes_3_4_io_outputA;
  wire       [7:0]    pes_3_4_io_outputB;
  wire       [25:0]   pes_3_4_io_outputC;
  wire       [7:0]    pes_3_5_io_outputA;
  wire       [7:0]    pes_3_5_io_outputB;
  wire       [25:0]   pes_3_5_io_outputC;
  wire       [7:0]    pes_3_6_io_outputA;
  wire       [7:0]    pes_3_6_io_outputB;
  wire       [25:0]   pes_3_6_io_outputC;
  wire       [7:0]    pes_3_7_io_outputA;
  wire       [7:0]    pes_3_7_io_outputB;
  wire       [25:0]   pes_3_7_io_outputC;
  wire       [7:0]    pes_3_8_io_outputA;
  wire       [7:0]    pes_3_8_io_outputB;
  wire       [25:0]   pes_3_8_io_outputC;
  wire       [7:0]    pes_3_9_io_outputA;
  wire       [7:0]    pes_3_9_io_outputB;
  wire       [25:0]   pes_3_9_io_outputC;
  wire       [7:0]    pes_3_10_io_outputA;
  wire       [7:0]    pes_3_10_io_outputB;
  wire       [25:0]   pes_3_10_io_outputC;
  wire       [7:0]    pes_3_11_io_outputA;
  wire       [7:0]    pes_3_11_io_outputB;
  wire       [25:0]   pes_3_11_io_outputC;
  wire       [7:0]    pes_3_12_io_outputA;
  wire       [7:0]    pes_3_12_io_outputB;
  wire       [25:0]   pes_3_12_io_outputC;
  wire       [7:0]    pes_3_13_io_outputA;
  wire       [7:0]    pes_3_13_io_outputB;
  wire       [25:0]   pes_3_13_io_outputC;
  wire       [7:0]    pes_3_14_io_outputA;
  wire       [7:0]    pes_3_14_io_outputB;
  wire       [25:0]   pes_3_14_io_outputC;
  wire       [7:0]    pes_3_15_io_outputB;
  wire       [25:0]   pes_3_15_io_outputC;
  wire       [7:0]    pes_4_0_io_outputA;
  wire       [7:0]    pes_4_0_io_outputB;
  wire       [25:0]   pes_4_0_io_outputC;
  wire       [7:0]    pes_4_1_io_outputA;
  wire       [7:0]    pes_4_1_io_outputB;
  wire       [25:0]   pes_4_1_io_outputC;
  wire       [7:0]    pes_4_2_io_outputA;
  wire       [7:0]    pes_4_2_io_outputB;
  wire       [25:0]   pes_4_2_io_outputC;
  wire       [7:0]    pes_4_3_io_outputA;
  wire       [7:0]    pes_4_3_io_outputB;
  wire       [25:0]   pes_4_3_io_outputC;
  wire       [7:0]    pes_4_4_io_outputA;
  wire       [7:0]    pes_4_4_io_outputB;
  wire       [25:0]   pes_4_4_io_outputC;
  wire       [7:0]    pes_4_5_io_outputA;
  wire       [7:0]    pes_4_5_io_outputB;
  wire       [25:0]   pes_4_5_io_outputC;
  wire       [7:0]    pes_4_6_io_outputA;
  wire       [7:0]    pes_4_6_io_outputB;
  wire       [25:0]   pes_4_6_io_outputC;
  wire       [7:0]    pes_4_7_io_outputA;
  wire       [7:0]    pes_4_7_io_outputB;
  wire       [25:0]   pes_4_7_io_outputC;
  wire       [7:0]    pes_4_8_io_outputA;
  wire       [7:0]    pes_4_8_io_outputB;
  wire       [25:0]   pes_4_8_io_outputC;
  wire       [7:0]    pes_4_9_io_outputA;
  wire       [7:0]    pes_4_9_io_outputB;
  wire       [25:0]   pes_4_9_io_outputC;
  wire       [7:0]    pes_4_10_io_outputA;
  wire       [7:0]    pes_4_10_io_outputB;
  wire       [25:0]   pes_4_10_io_outputC;
  wire       [7:0]    pes_4_11_io_outputA;
  wire       [7:0]    pes_4_11_io_outputB;
  wire       [25:0]   pes_4_11_io_outputC;
  wire       [7:0]    pes_4_12_io_outputA;
  wire       [7:0]    pes_4_12_io_outputB;
  wire       [25:0]   pes_4_12_io_outputC;
  wire       [7:0]    pes_4_13_io_outputA;
  wire       [7:0]    pes_4_13_io_outputB;
  wire       [25:0]   pes_4_13_io_outputC;
  wire       [7:0]    pes_4_14_io_outputA;
  wire       [7:0]    pes_4_14_io_outputB;
  wire       [25:0]   pes_4_14_io_outputC;
  wire       [7:0]    pes_4_15_io_outputB;
  wire       [25:0]   pes_4_15_io_outputC;
  wire       [7:0]    pes_5_0_io_outputA;
  wire       [7:0]    pes_5_0_io_outputB;
  wire       [25:0]   pes_5_0_io_outputC;
  wire       [7:0]    pes_5_1_io_outputA;
  wire       [7:0]    pes_5_1_io_outputB;
  wire       [25:0]   pes_5_1_io_outputC;
  wire       [7:0]    pes_5_2_io_outputA;
  wire       [7:0]    pes_5_2_io_outputB;
  wire       [25:0]   pes_5_2_io_outputC;
  wire       [7:0]    pes_5_3_io_outputA;
  wire       [7:0]    pes_5_3_io_outputB;
  wire       [25:0]   pes_5_3_io_outputC;
  wire       [7:0]    pes_5_4_io_outputA;
  wire       [7:0]    pes_5_4_io_outputB;
  wire       [25:0]   pes_5_4_io_outputC;
  wire       [7:0]    pes_5_5_io_outputA;
  wire       [7:0]    pes_5_5_io_outputB;
  wire       [25:0]   pes_5_5_io_outputC;
  wire       [7:0]    pes_5_6_io_outputA;
  wire       [7:0]    pes_5_6_io_outputB;
  wire       [25:0]   pes_5_6_io_outputC;
  wire       [7:0]    pes_5_7_io_outputA;
  wire       [7:0]    pes_5_7_io_outputB;
  wire       [25:0]   pes_5_7_io_outputC;
  wire       [7:0]    pes_5_8_io_outputA;
  wire       [7:0]    pes_5_8_io_outputB;
  wire       [25:0]   pes_5_8_io_outputC;
  wire       [7:0]    pes_5_9_io_outputA;
  wire       [7:0]    pes_5_9_io_outputB;
  wire       [25:0]   pes_5_9_io_outputC;
  wire       [7:0]    pes_5_10_io_outputA;
  wire       [7:0]    pes_5_10_io_outputB;
  wire       [25:0]   pes_5_10_io_outputC;
  wire       [7:0]    pes_5_11_io_outputA;
  wire       [7:0]    pes_5_11_io_outputB;
  wire       [25:0]   pes_5_11_io_outputC;
  wire       [7:0]    pes_5_12_io_outputA;
  wire       [7:0]    pes_5_12_io_outputB;
  wire       [25:0]   pes_5_12_io_outputC;
  wire       [7:0]    pes_5_13_io_outputA;
  wire       [7:0]    pes_5_13_io_outputB;
  wire       [25:0]   pes_5_13_io_outputC;
  wire       [7:0]    pes_5_14_io_outputA;
  wire       [7:0]    pes_5_14_io_outputB;
  wire       [25:0]   pes_5_14_io_outputC;
  wire       [7:0]    pes_5_15_io_outputB;
  wire       [25:0]   pes_5_15_io_outputC;
  wire       [7:0]    pes_6_0_io_outputA;
  wire       [7:0]    pes_6_0_io_outputB;
  wire       [25:0]   pes_6_0_io_outputC;
  wire       [7:0]    pes_6_1_io_outputA;
  wire       [7:0]    pes_6_1_io_outputB;
  wire       [25:0]   pes_6_1_io_outputC;
  wire       [7:0]    pes_6_2_io_outputA;
  wire       [7:0]    pes_6_2_io_outputB;
  wire       [25:0]   pes_6_2_io_outputC;
  wire       [7:0]    pes_6_3_io_outputA;
  wire       [7:0]    pes_6_3_io_outputB;
  wire       [25:0]   pes_6_3_io_outputC;
  wire       [7:0]    pes_6_4_io_outputA;
  wire       [7:0]    pes_6_4_io_outputB;
  wire       [25:0]   pes_6_4_io_outputC;
  wire       [7:0]    pes_6_5_io_outputA;
  wire       [7:0]    pes_6_5_io_outputB;
  wire       [25:0]   pes_6_5_io_outputC;
  wire       [7:0]    pes_6_6_io_outputA;
  wire       [7:0]    pes_6_6_io_outputB;
  wire       [25:0]   pes_6_6_io_outputC;
  wire       [7:0]    pes_6_7_io_outputA;
  wire       [7:0]    pes_6_7_io_outputB;
  wire       [25:0]   pes_6_7_io_outputC;
  wire       [7:0]    pes_6_8_io_outputA;
  wire       [7:0]    pes_6_8_io_outputB;
  wire       [25:0]   pes_6_8_io_outputC;
  wire       [7:0]    pes_6_9_io_outputA;
  wire       [7:0]    pes_6_9_io_outputB;
  wire       [25:0]   pes_6_9_io_outputC;
  wire       [7:0]    pes_6_10_io_outputA;
  wire       [7:0]    pes_6_10_io_outputB;
  wire       [25:0]   pes_6_10_io_outputC;
  wire       [7:0]    pes_6_11_io_outputA;
  wire       [7:0]    pes_6_11_io_outputB;
  wire       [25:0]   pes_6_11_io_outputC;
  wire       [7:0]    pes_6_12_io_outputA;
  wire       [7:0]    pes_6_12_io_outputB;
  wire       [25:0]   pes_6_12_io_outputC;
  wire       [7:0]    pes_6_13_io_outputA;
  wire       [7:0]    pes_6_13_io_outputB;
  wire       [25:0]   pes_6_13_io_outputC;
  wire       [7:0]    pes_6_14_io_outputA;
  wire       [7:0]    pes_6_14_io_outputB;
  wire       [25:0]   pes_6_14_io_outputC;
  wire       [7:0]    pes_6_15_io_outputB;
  wire       [25:0]   pes_6_15_io_outputC;
  wire       [7:0]    pes_7_0_io_outputA;
  wire       [7:0]    pes_7_0_io_outputB;
  wire       [25:0]   pes_7_0_io_outputC;
  wire       [7:0]    pes_7_1_io_outputA;
  wire       [7:0]    pes_7_1_io_outputB;
  wire       [25:0]   pes_7_1_io_outputC;
  wire       [7:0]    pes_7_2_io_outputA;
  wire       [7:0]    pes_7_2_io_outputB;
  wire       [25:0]   pes_7_2_io_outputC;
  wire       [7:0]    pes_7_3_io_outputA;
  wire       [7:0]    pes_7_3_io_outputB;
  wire       [25:0]   pes_7_3_io_outputC;
  wire       [7:0]    pes_7_4_io_outputA;
  wire       [7:0]    pes_7_4_io_outputB;
  wire       [25:0]   pes_7_4_io_outputC;
  wire       [7:0]    pes_7_5_io_outputA;
  wire       [7:0]    pes_7_5_io_outputB;
  wire       [25:0]   pes_7_5_io_outputC;
  wire       [7:0]    pes_7_6_io_outputA;
  wire       [7:0]    pes_7_6_io_outputB;
  wire       [25:0]   pes_7_6_io_outputC;
  wire       [7:0]    pes_7_7_io_outputA;
  wire       [7:0]    pes_7_7_io_outputB;
  wire       [25:0]   pes_7_7_io_outputC;
  wire       [7:0]    pes_7_8_io_outputA;
  wire       [7:0]    pes_7_8_io_outputB;
  wire       [25:0]   pes_7_8_io_outputC;
  wire       [7:0]    pes_7_9_io_outputA;
  wire       [7:0]    pes_7_9_io_outputB;
  wire       [25:0]   pes_7_9_io_outputC;
  wire       [7:0]    pes_7_10_io_outputA;
  wire       [7:0]    pes_7_10_io_outputB;
  wire       [25:0]   pes_7_10_io_outputC;
  wire       [7:0]    pes_7_11_io_outputA;
  wire       [7:0]    pes_7_11_io_outputB;
  wire       [25:0]   pes_7_11_io_outputC;
  wire       [7:0]    pes_7_12_io_outputA;
  wire       [7:0]    pes_7_12_io_outputB;
  wire       [25:0]   pes_7_12_io_outputC;
  wire       [7:0]    pes_7_13_io_outputA;
  wire       [7:0]    pes_7_13_io_outputB;
  wire       [25:0]   pes_7_13_io_outputC;
  wire       [7:0]    pes_7_14_io_outputA;
  wire       [7:0]    pes_7_14_io_outputB;
  wire       [25:0]   pes_7_14_io_outputC;
  wire       [7:0]    pes_7_15_io_outputB;
  wire       [25:0]   pes_7_15_io_outputC;
  wire       [7:0]    pes_8_0_io_outputA;
  wire       [7:0]    pes_8_0_io_outputB;
  wire       [25:0]   pes_8_0_io_outputC;
  wire       [7:0]    pes_8_1_io_outputA;
  wire       [7:0]    pes_8_1_io_outputB;
  wire       [25:0]   pes_8_1_io_outputC;
  wire       [7:0]    pes_8_2_io_outputA;
  wire       [7:0]    pes_8_2_io_outputB;
  wire       [25:0]   pes_8_2_io_outputC;
  wire       [7:0]    pes_8_3_io_outputA;
  wire       [7:0]    pes_8_3_io_outputB;
  wire       [25:0]   pes_8_3_io_outputC;
  wire       [7:0]    pes_8_4_io_outputA;
  wire       [7:0]    pes_8_4_io_outputB;
  wire       [25:0]   pes_8_4_io_outputC;
  wire       [7:0]    pes_8_5_io_outputA;
  wire       [7:0]    pes_8_5_io_outputB;
  wire       [25:0]   pes_8_5_io_outputC;
  wire       [7:0]    pes_8_6_io_outputA;
  wire       [7:0]    pes_8_6_io_outputB;
  wire       [25:0]   pes_8_6_io_outputC;
  wire       [7:0]    pes_8_7_io_outputA;
  wire       [7:0]    pes_8_7_io_outputB;
  wire       [25:0]   pes_8_7_io_outputC;
  wire       [7:0]    pes_8_8_io_outputA;
  wire       [7:0]    pes_8_8_io_outputB;
  wire       [25:0]   pes_8_8_io_outputC;
  wire       [7:0]    pes_8_9_io_outputA;
  wire       [7:0]    pes_8_9_io_outputB;
  wire       [25:0]   pes_8_9_io_outputC;
  wire       [7:0]    pes_8_10_io_outputA;
  wire       [7:0]    pes_8_10_io_outputB;
  wire       [25:0]   pes_8_10_io_outputC;
  wire       [7:0]    pes_8_11_io_outputA;
  wire       [7:0]    pes_8_11_io_outputB;
  wire       [25:0]   pes_8_11_io_outputC;
  wire       [7:0]    pes_8_12_io_outputA;
  wire       [7:0]    pes_8_12_io_outputB;
  wire       [25:0]   pes_8_12_io_outputC;
  wire       [7:0]    pes_8_13_io_outputA;
  wire       [7:0]    pes_8_13_io_outputB;
  wire       [25:0]   pes_8_13_io_outputC;
  wire       [7:0]    pes_8_14_io_outputA;
  wire       [7:0]    pes_8_14_io_outputB;
  wire       [25:0]   pes_8_14_io_outputC;
  wire       [7:0]    pes_8_15_io_outputB;
  wire       [25:0]   pes_8_15_io_outputC;
  wire       [7:0]    pes_9_0_io_outputA;
  wire       [7:0]    pes_9_0_io_outputB;
  wire       [25:0]   pes_9_0_io_outputC;
  wire       [7:0]    pes_9_1_io_outputA;
  wire       [7:0]    pes_9_1_io_outputB;
  wire       [25:0]   pes_9_1_io_outputC;
  wire       [7:0]    pes_9_2_io_outputA;
  wire       [7:0]    pes_9_2_io_outputB;
  wire       [25:0]   pes_9_2_io_outputC;
  wire       [7:0]    pes_9_3_io_outputA;
  wire       [7:0]    pes_9_3_io_outputB;
  wire       [25:0]   pes_9_3_io_outputC;
  wire       [7:0]    pes_9_4_io_outputA;
  wire       [7:0]    pes_9_4_io_outputB;
  wire       [25:0]   pes_9_4_io_outputC;
  wire       [7:0]    pes_9_5_io_outputA;
  wire       [7:0]    pes_9_5_io_outputB;
  wire       [25:0]   pes_9_5_io_outputC;
  wire       [7:0]    pes_9_6_io_outputA;
  wire       [7:0]    pes_9_6_io_outputB;
  wire       [25:0]   pes_9_6_io_outputC;
  wire       [7:0]    pes_9_7_io_outputA;
  wire       [7:0]    pes_9_7_io_outputB;
  wire       [25:0]   pes_9_7_io_outputC;
  wire       [7:0]    pes_9_8_io_outputA;
  wire       [7:0]    pes_9_8_io_outputB;
  wire       [25:0]   pes_9_8_io_outputC;
  wire       [7:0]    pes_9_9_io_outputA;
  wire       [7:0]    pes_9_9_io_outputB;
  wire       [25:0]   pes_9_9_io_outputC;
  wire       [7:0]    pes_9_10_io_outputA;
  wire       [7:0]    pes_9_10_io_outputB;
  wire       [25:0]   pes_9_10_io_outputC;
  wire       [7:0]    pes_9_11_io_outputA;
  wire       [7:0]    pes_9_11_io_outputB;
  wire       [25:0]   pes_9_11_io_outputC;
  wire       [7:0]    pes_9_12_io_outputA;
  wire       [7:0]    pes_9_12_io_outputB;
  wire       [25:0]   pes_9_12_io_outputC;
  wire       [7:0]    pes_9_13_io_outputA;
  wire       [7:0]    pes_9_13_io_outputB;
  wire       [25:0]   pes_9_13_io_outputC;
  wire       [7:0]    pes_9_14_io_outputA;
  wire       [7:0]    pes_9_14_io_outputB;
  wire       [25:0]   pes_9_14_io_outputC;
  wire       [7:0]    pes_9_15_io_outputB;
  wire       [25:0]   pes_9_15_io_outputC;
  wire       [7:0]    pes_10_0_io_outputA;
  wire       [7:0]    pes_10_0_io_outputB;
  wire       [25:0]   pes_10_0_io_outputC;
  wire       [7:0]    pes_10_1_io_outputA;
  wire       [7:0]    pes_10_1_io_outputB;
  wire       [25:0]   pes_10_1_io_outputC;
  wire       [7:0]    pes_10_2_io_outputA;
  wire       [7:0]    pes_10_2_io_outputB;
  wire       [25:0]   pes_10_2_io_outputC;
  wire       [7:0]    pes_10_3_io_outputA;
  wire       [7:0]    pes_10_3_io_outputB;
  wire       [25:0]   pes_10_3_io_outputC;
  wire       [7:0]    pes_10_4_io_outputA;
  wire       [7:0]    pes_10_4_io_outputB;
  wire       [25:0]   pes_10_4_io_outputC;
  wire       [7:0]    pes_10_5_io_outputA;
  wire       [7:0]    pes_10_5_io_outputB;
  wire       [25:0]   pes_10_5_io_outputC;
  wire       [7:0]    pes_10_6_io_outputA;
  wire       [7:0]    pes_10_6_io_outputB;
  wire       [25:0]   pes_10_6_io_outputC;
  wire       [7:0]    pes_10_7_io_outputA;
  wire       [7:0]    pes_10_7_io_outputB;
  wire       [25:0]   pes_10_7_io_outputC;
  wire       [7:0]    pes_10_8_io_outputA;
  wire       [7:0]    pes_10_8_io_outputB;
  wire       [25:0]   pes_10_8_io_outputC;
  wire       [7:0]    pes_10_9_io_outputA;
  wire       [7:0]    pes_10_9_io_outputB;
  wire       [25:0]   pes_10_9_io_outputC;
  wire       [7:0]    pes_10_10_io_outputA;
  wire       [7:0]    pes_10_10_io_outputB;
  wire       [25:0]   pes_10_10_io_outputC;
  wire       [7:0]    pes_10_11_io_outputA;
  wire       [7:0]    pes_10_11_io_outputB;
  wire       [25:0]   pes_10_11_io_outputC;
  wire       [7:0]    pes_10_12_io_outputA;
  wire       [7:0]    pes_10_12_io_outputB;
  wire       [25:0]   pes_10_12_io_outputC;
  wire       [7:0]    pes_10_13_io_outputA;
  wire       [7:0]    pes_10_13_io_outputB;
  wire       [25:0]   pes_10_13_io_outputC;
  wire       [7:0]    pes_10_14_io_outputA;
  wire       [7:0]    pes_10_14_io_outputB;
  wire       [25:0]   pes_10_14_io_outputC;
  wire       [7:0]    pes_10_15_io_outputB;
  wire       [25:0]   pes_10_15_io_outputC;
  wire       [7:0]    pes_11_0_io_outputA;
  wire       [7:0]    pes_11_0_io_outputB;
  wire       [25:0]   pes_11_0_io_outputC;
  wire       [7:0]    pes_11_1_io_outputA;
  wire       [7:0]    pes_11_1_io_outputB;
  wire       [25:0]   pes_11_1_io_outputC;
  wire       [7:0]    pes_11_2_io_outputA;
  wire       [7:0]    pes_11_2_io_outputB;
  wire       [25:0]   pes_11_2_io_outputC;
  wire       [7:0]    pes_11_3_io_outputA;
  wire       [7:0]    pes_11_3_io_outputB;
  wire       [25:0]   pes_11_3_io_outputC;
  wire       [7:0]    pes_11_4_io_outputA;
  wire       [7:0]    pes_11_4_io_outputB;
  wire       [25:0]   pes_11_4_io_outputC;
  wire       [7:0]    pes_11_5_io_outputA;
  wire       [7:0]    pes_11_5_io_outputB;
  wire       [25:0]   pes_11_5_io_outputC;
  wire       [7:0]    pes_11_6_io_outputA;
  wire       [7:0]    pes_11_6_io_outputB;
  wire       [25:0]   pes_11_6_io_outputC;
  wire       [7:0]    pes_11_7_io_outputA;
  wire       [7:0]    pes_11_7_io_outputB;
  wire       [25:0]   pes_11_7_io_outputC;
  wire       [7:0]    pes_11_8_io_outputA;
  wire       [7:0]    pes_11_8_io_outputB;
  wire       [25:0]   pes_11_8_io_outputC;
  wire       [7:0]    pes_11_9_io_outputA;
  wire       [7:0]    pes_11_9_io_outputB;
  wire       [25:0]   pes_11_9_io_outputC;
  wire       [7:0]    pes_11_10_io_outputA;
  wire       [7:0]    pes_11_10_io_outputB;
  wire       [25:0]   pes_11_10_io_outputC;
  wire       [7:0]    pes_11_11_io_outputA;
  wire       [7:0]    pes_11_11_io_outputB;
  wire       [25:0]   pes_11_11_io_outputC;
  wire       [7:0]    pes_11_12_io_outputA;
  wire       [7:0]    pes_11_12_io_outputB;
  wire       [25:0]   pes_11_12_io_outputC;
  wire       [7:0]    pes_11_13_io_outputA;
  wire       [7:0]    pes_11_13_io_outputB;
  wire       [25:0]   pes_11_13_io_outputC;
  wire       [7:0]    pes_11_14_io_outputA;
  wire       [7:0]    pes_11_14_io_outputB;
  wire       [25:0]   pes_11_14_io_outputC;
  wire       [7:0]    pes_11_15_io_outputB;
  wire       [25:0]   pes_11_15_io_outputC;
  wire       [7:0]    pes_12_0_io_outputA;
  wire       [7:0]    pes_12_0_io_outputB;
  wire       [25:0]   pes_12_0_io_outputC;
  wire       [7:0]    pes_12_1_io_outputA;
  wire       [7:0]    pes_12_1_io_outputB;
  wire       [25:0]   pes_12_1_io_outputC;
  wire       [7:0]    pes_12_2_io_outputA;
  wire       [7:0]    pes_12_2_io_outputB;
  wire       [25:0]   pes_12_2_io_outputC;
  wire       [7:0]    pes_12_3_io_outputA;
  wire       [7:0]    pes_12_3_io_outputB;
  wire       [25:0]   pes_12_3_io_outputC;
  wire       [7:0]    pes_12_4_io_outputA;
  wire       [7:0]    pes_12_4_io_outputB;
  wire       [25:0]   pes_12_4_io_outputC;
  wire       [7:0]    pes_12_5_io_outputA;
  wire       [7:0]    pes_12_5_io_outputB;
  wire       [25:0]   pes_12_5_io_outputC;
  wire       [7:0]    pes_12_6_io_outputA;
  wire       [7:0]    pes_12_6_io_outputB;
  wire       [25:0]   pes_12_6_io_outputC;
  wire       [7:0]    pes_12_7_io_outputA;
  wire       [7:0]    pes_12_7_io_outputB;
  wire       [25:0]   pes_12_7_io_outputC;
  wire       [7:0]    pes_12_8_io_outputA;
  wire       [7:0]    pes_12_8_io_outputB;
  wire       [25:0]   pes_12_8_io_outputC;
  wire       [7:0]    pes_12_9_io_outputA;
  wire       [7:0]    pes_12_9_io_outputB;
  wire       [25:0]   pes_12_9_io_outputC;
  wire       [7:0]    pes_12_10_io_outputA;
  wire       [7:0]    pes_12_10_io_outputB;
  wire       [25:0]   pes_12_10_io_outputC;
  wire       [7:0]    pes_12_11_io_outputA;
  wire       [7:0]    pes_12_11_io_outputB;
  wire       [25:0]   pes_12_11_io_outputC;
  wire       [7:0]    pes_12_12_io_outputA;
  wire       [7:0]    pes_12_12_io_outputB;
  wire       [25:0]   pes_12_12_io_outputC;
  wire       [7:0]    pes_12_13_io_outputA;
  wire       [7:0]    pes_12_13_io_outputB;
  wire       [25:0]   pes_12_13_io_outputC;
  wire       [7:0]    pes_12_14_io_outputA;
  wire       [7:0]    pes_12_14_io_outputB;
  wire       [25:0]   pes_12_14_io_outputC;
  wire       [7:0]    pes_12_15_io_outputB;
  wire       [25:0]   pes_12_15_io_outputC;
  wire       [7:0]    pes_13_0_io_outputA;
  wire       [7:0]    pes_13_0_io_outputB;
  wire       [25:0]   pes_13_0_io_outputC;
  wire       [7:0]    pes_13_1_io_outputA;
  wire       [7:0]    pes_13_1_io_outputB;
  wire       [25:0]   pes_13_1_io_outputC;
  wire       [7:0]    pes_13_2_io_outputA;
  wire       [7:0]    pes_13_2_io_outputB;
  wire       [25:0]   pes_13_2_io_outputC;
  wire       [7:0]    pes_13_3_io_outputA;
  wire       [7:0]    pes_13_3_io_outputB;
  wire       [25:0]   pes_13_3_io_outputC;
  wire       [7:0]    pes_13_4_io_outputA;
  wire       [7:0]    pes_13_4_io_outputB;
  wire       [25:0]   pes_13_4_io_outputC;
  wire       [7:0]    pes_13_5_io_outputA;
  wire       [7:0]    pes_13_5_io_outputB;
  wire       [25:0]   pes_13_5_io_outputC;
  wire       [7:0]    pes_13_6_io_outputA;
  wire       [7:0]    pes_13_6_io_outputB;
  wire       [25:0]   pes_13_6_io_outputC;
  wire       [7:0]    pes_13_7_io_outputA;
  wire       [7:0]    pes_13_7_io_outputB;
  wire       [25:0]   pes_13_7_io_outputC;
  wire       [7:0]    pes_13_8_io_outputA;
  wire       [7:0]    pes_13_8_io_outputB;
  wire       [25:0]   pes_13_8_io_outputC;
  wire       [7:0]    pes_13_9_io_outputA;
  wire       [7:0]    pes_13_9_io_outputB;
  wire       [25:0]   pes_13_9_io_outputC;
  wire       [7:0]    pes_13_10_io_outputA;
  wire       [7:0]    pes_13_10_io_outputB;
  wire       [25:0]   pes_13_10_io_outputC;
  wire       [7:0]    pes_13_11_io_outputA;
  wire       [7:0]    pes_13_11_io_outputB;
  wire       [25:0]   pes_13_11_io_outputC;
  wire       [7:0]    pes_13_12_io_outputA;
  wire       [7:0]    pes_13_12_io_outputB;
  wire       [25:0]   pes_13_12_io_outputC;
  wire       [7:0]    pes_13_13_io_outputA;
  wire       [7:0]    pes_13_13_io_outputB;
  wire       [25:0]   pes_13_13_io_outputC;
  wire       [7:0]    pes_13_14_io_outputA;
  wire       [7:0]    pes_13_14_io_outputB;
  wire       [25:0]   pes_13_14_io_outputC;
  wire       [7:0]    pes_13_15_io_outputB;
  wire       [25:0]   pes_13_15_io_outputC;
  wire       [7:0]    pes_14_0_io_outputA;
  wire       [7:0]    pes_14_0_io_outputB;
  wire       [25:0]   pes_14_0_io_outputC;
  wire       [7:0]    pes_14_1_io_outputA;
  wire       [7:0]    pes_14_1_io_outputB;
  wire       [25:0]   pes_14_1_io_outputC;
  wire       [7:0]    pes_14_2_io_outputA;
  wire       [7:0]    pes_14_2_io_outputB;
  wire       [25:0]   pes_14_2_io_outputC;
  wire       [7:0]    pes_14_3_io_outputA;
  wire       [7:0]    pes_14_3_io_outputB;
  wire       [25:0]   pes_14_3_io_outputC;
  wire       [7:0]    pes_14_4_io_outputA;
  wire       [7:0]    pes_14_4_io_outputB;
  wire       [25:0]   pes_14_4_io_outputC;
  wire       [7:0]    pes_14_5_io_outputA;
  wire       [7:0]    pes_14_5_io_outputB;
  wire       [25:0]   pes_14_5_io_outputC;
  wire       [7:0]    pes_14_6_io_outputA;
  wire       [7:0]    pes_14_6_io_outputB;
  wire       [25:0]   pes_14_6_io_outputC;
  wire       [7:0]    pes_14_7_io_outputA;
  wire       [7:0]    pes_14_7_io_outputB;
  wire       [25:0]   pes_14_7_io_outputC;
  wire       [7:0]    pes_14_8_io_outputA;
  wire       [7:0]    pes_14_8_io_outputB;
  wire       [25:0]   pes_14_8_io_outputC;
  wire       [7:0]    pes_14_9_io_outputA;
  wire       [7:0]    pes_14_9_io_outputB;
  wire       [25:0]   pes_14_9_io_outputC;
  wire       [7:0]    pes_14_10_io_outputA;
  wire       [7:0]    pes_14_10_io_outputB;
  wire       [25:0]   pes_14_10_io_outputC;
  wire       [7:0]    pes_14_11_io_outputA;
  wire       [7:0]    pes_14_11_io_outputB;
  wire       [25:0]   pes_14_11_io_outputC;
  wire       [7:0]    pes_14_12_io_outputA;
  wire       [7:0]    pes_14_12_io_outputB;
  wire       [25:0]   pes_14_12_io_outputC;
  wire       [7:0]    pes_14_13_io_outputA;
  wire       [7:0]    pes_14_13_io_outputB;
  wire       [25:0]   pes_14_13_io_outputC;
  wire       [7:0]    pes_14_14_io_outputA;
  wire       [7:0]    pes_14_14_io_outputB;
  wire       [25:0]   pes_14_14_io_outputC;
  wire       [7:0]    pes_14_15_io_outputB;
  wire       [25:0]   pes_14_15_io_outputC;
  wire       [7:0]    pes_15_0_io_outputA;
  wire       [25:0]   pes_15_0_io_outputC;
  wire       [7:0]    pes_15_1_io_outputA;
  wire       [25:0]   pes_15_1_io_outputC;
  wire       [7:0]    pes_15_2_io_outputA;
  wire       [25:0]   pes_15_2_io_outputC;
  wire       [7:0]    pes_15_3_io_outputA;
  wire       [25:0]   pes_15_3_io_outputC;
  wire       [7:0]    pes_15_4_io_outputA;
  wire       [25:0]   pes_15_4_io_outputC;
  wire       [7:0]    pes_15_5_io_outputA;
  wire       [25:0]   pes_15_5_io_outputC;
  wire       [7:0]    pes_15_6_io_outputA;
  wire       [25:0]   pes_15_6_io_outputC;
  wire       [7:0]    pes_15_7_io_outputA;
  wire       [25:0]   pes_15_7_io_outputC;
  wire       [7:0]    pes_15_8_io_outputA;
  wire       [25:0]   pes_15_8_io_outputC;
  wire       [7:0]    pes_15_9_io_outputA;
  wire       [25:0]   pes_15_9_io_outputC;
  wire       [7:0]    pes_15_10_io_outputA;
  wire       [25:0]   pes_15_10_io_outputC;
  wire       [7:0]    pes_15_11_io_outputA;
  wire       [25:0]   pes_15_11_io_outputC;
  wire       [7:0]    pes_15_12_io_outputA;
  wire       [25:0]   pes_15_12_io_outputC;
  wire       [7:0]    pes_15_13_io_outputA;
  wire       [25:0]   pes_15_13_io_outputC;
  wire       [7:0]    pes_15_14_io_outputA;
  wire       [25:0]   pes_15_14_io_outputC;
  wire       [25:0]   pes_15_15_io_outputC;
  wire       [7:0]    skewBuffer_io_output_0;
  wire       [7:0]    skewBuffer_io_output_1;
  wire       [7:0]    skewBuffer_io_output_2;
  wire       [7:0]    skewBuffer_io_output_3;
  wire       [7:0]    skewBuffer_io_output_4;
  wire       [7:0]    skewBuffer_io_output_5;
  wire       [7:0]    skewBuffer_io_output_6;
  wire       [7:0]    skewBuffer_io_output_7;
  wire       [7:0]    skewBuffer_io_output_8;
  wire       [7:0]    skewBuffer_io_output_9;
  wire       [7:0]    skewBuffer_io_output_10;
  wire       [7:0]    skewBuffer_io_output_11;
  wire       [7:0]    skewBuffer_io_output_12;
  wire       [7:0]    skewBuffer_io_output_13;
  wire       [7:0]    skewBuffer_io_output_14;
  wire       [7:0]    skewBuffer_io_output_15;
  wire       [7:0]    skewBuffer_1_io_output_0;
  wire       [7:0]    skewBuffer_1_io_output_1;
  wire       [7:0]    skewBuffer_1_io_output_2;
  wire       [7:0]    skewBuffer_1_io_output_3;
  wire       [7:0]    skewBuffer_1_io_output_4;
  wire       [7:0]    skewBuffer_1_io_output_5;
  wire       [7:0]    skewBuffer_1_io_output_6;
  wire       [7:0]    skewBuffer_1_io_output_7;
  wire       [7:0]    skewBuffer_1_io_output_8;
  wire       [7:0]    skewBuffer_1_io_output_9;
  wire       [7:0]    skewBuffer_1_io_output_10;
  wire       [7:0]    skewBuffer_1_io_output_11;
  wire       [7:0]    skewBuffer_1_io_output_12;
  wire       [7:0]    skewBuffer_1_io_output_13;
  wire       [7:0]    skewBuffer_1_io_output_14;
  wire       [7:0]    skewBuffer_1_io_output_15;
  wire       [25:0]   deskewBufferReuseC_io_output_0;
  wire       [25:0]   deskewBufferReuseC_io_output_1;
  wire       [25:0]   deskewBufferReuseC_io_output_2;
  wire       [25:0]   deskewBufferReuseC_io_output_3;
  wire       [25:0]   deskewBufferReuseC_io_output_4;
  wire       [25:0]   deskewBufferReuseC_io_output_5;
  wire       [25:0]   deskewBufferReuseC_io_output_6;
  wire       [25:0]   deskewBufferReuseC_io_output_7;
  wire       [25:0]   deskewBufferReuseC_io_output_8;
  wire       [25:0]   deskewBufferReuseC_io_output_9;
  wire       [25:0]   deskewBufferReuseC_io_output_10;
  wire       [25:0]   deskewBufferReuseC_io_output_11;
  wire       [25:0]   deskewBufferReuseC_io_output_12;
  wire       [25:0]   deskewBufferReuseC_io_output_13;
  wire       [25:0]   deskewBufferReuseC_io_output_14;
  wire       [25:0]   deskewBufferReuseC_io_output_15;
  wire       [25:0]   deskewBufferReuseC_io_output_16;
  wire       [25:0]   deskewBufferReuseC_io_output_17;
  wire       [25:0]   deskewBufferReuseC_io_output_18;
  wire       [25:0]   deskewBufferReuseC_io_output_19;
  wire       [25:0]   deskewBufferReuseC_io_output_20;
  wire       [25:0]   deskewBufferReuseC_io_output_21;
  wire       [25:0]   deskewBufferReuseC_io_output_22;
  wire       [25:0]   deskewBufferReuseC_io_output_23;
  wire       [25:0]   deskewBufferReuseC_io_output_24;
  wire       [25:0]   deskewBufferReuseC_io_output_25;
  wire       [25:0]   deskewBufferReuseC_io_output_26;
  wire       [25:0]   deskewBufferReuseC_io_output_27;
  wire       [25:0]   deskewBufferReuseC_io_output_28;
  wire       [25:0]   deskewBufferReuseC_io_output_29;
  wire       [25:0]   deskewBufferReuseC_io_output_30;

  ProcessingElement pes_0_0 (
    .io_inputA               (skewBuffer_io_output_0[7:0]  ), //i
    .io_inputB               (skewBuffer_1_io_output_0[7:0]), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_0_0  ), //i
    .io_resetPartialC        (io_resetPartialC_0_0         ), //i
    .io_outputA              (pes_0_0_io_outputA[7:0]      ), //o
    .io_outputB              (pes_0_0_io_outputB[7:0]      ), //o
    .io_outputC              (pes_0_0_io_outputC[25:0]     ), //o
    .clk                     (clk                          ), //i
    .reset                   (reset                        )  //i
  );
  ProcessingElement pes_0_1 (
    .io_inputA               (pes_0_0_io_outputA[7:0]      ), //i
    .io_inputB               (skewBuffer_1_io_output_1[7:0]), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_0_1  ), //i
    .io_resetPartialC        (io_resetPartialC_0_1         ), //i
    .io_outputA              (pes_0_1_io_outputA[7:0]      ), //o
    .io_outputB              (pes_0_1_io_outputB[7:0]      ), //o
    .io_outputC              (pes_0_1_io_outputC[25:0]     ), //o
    .clk                     (clk                          ), //i
    .reset                   (reset                        )  //i
  );
  ProcessingElement pes_0_2 (
    .io_inputA               (pes_0_1_io_outputA[7:0]      ), //i
    .io_inputB               (skewBuffer_1_io_output_2[7:0]), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_0_2  ), //i
    .io_resetPartialC        (io_resetPartialC_0_2         ), //i
    .io_outputA              (pes_0_2_io_outputA[7:0]      ), //o
    .io_outputB              (pes_0_2_io_outputB[7:0]      ), //o
    .io_outputC              (pes_0_2_io_outputC[25:0]     ), //o
    .clk                     (clk                          ), //i
    .reset                   (reset                        )  //i
  );
  ProcessingElement pes_0_3 (
    .io_inputA               (pes_0_2_io_outputA[7:0]      ), //i
    .io_inputB               (skewBuffer_1_io_output_3[7:0]), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_0_3  ), //i
    .io_resetPartialC        (io_resetPartialC_0_3         ), //i
    .io_outputA              (pes_0_3_io_outputA[7:0]      ), //o
    .io_outputB              (pes_0_3_io_outputB[7:0]      ), //o
    .io_outputC              (pes_0_3_io_outputC[25:0]     ), //o
    .clk                     (clk                          ), //i
    .reset                   (reset                        )  //i
  );
  ProcessingElement pes_0_4 (
    .io_inputA               (pes_0_3_io_outputA[7:0]      ), //i
    .io_inputB               (skewBuffer_1_io_output_4[7:0]), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_0_4  ), //i
    .io_resetPartialC        (io_resetPartialC_0_4         ), //i
    .io_outputA              (pes_0_4_io_outputA[7:0]      ), //o
    .io_outputB              (pes_0_4_io_outputB[7:0]      ), //o
    .io_outputC              (pes_0_4_io_outputC[25:0]     ), //o
    .clk                     (clk                          ), //i
    .reset                   (reset                        )  //i
  );
  ProcessingElement pes_0_5 (
    .io_inputA               (pes_0_4_io_outputA[7:0]      ), //i
    .io_inputB               (skewBuffer_1_io_output_5[7:0]), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_0_5  ), //i
    .io_resetPartialC        (io_resetPartialC_0_5         ), //i
    .io_outputA              (pes_0_5_io_outputA[7:0]      ), //o
    .io_outputB              (pes_0_5_io_outputB[7:0]      ), //o
    .io_outputC              (pes_0_5_io_outputC[25:0]     ), //o
    .clk                     (clk                          ), //i
    .reset                   (reset                        )  //i
  );
  ProcessingElement pes_0_6 (
    .io_inputA               (pes_0_5_io_outputA[7:0]      ), //i
    .io_inputB               (skewBuffer_1_io_output_6[7:0]), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_0_6  ), //i
    .io_resetPartialC        (io_resetPartialC_0_6         ), //i
    .io_outputA              (pes_0_6_io_outputA[7:0]      ), //o
    .io_outputB              (pes_0_6_io_outputB[7:0]      ), //o
    .io_outputC              (pes_0_6_io_outputC[25:0]     ), //o
    .clk                     (clk                          ), //i
    .reset                   (reset                        )  //i
  );
  ProcessingElement pes_0_7 (
    .io_inputA               (pes_0_6_io_outputA[7:0]      ), //i
    .io_inputB               (skewBuffer_1_io_output_7[7:0]), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_0_7  ), //i
    .io_resetPartialC        (io_resetPartialC_0_7         ), //i
    .io_outputA              (pes_0_7_io_outputA[7:0]      ), //o
    .io_outputB              (pes_0_7_io_outputB[7:0]      ), //o
    .io_outputC              (pes_0_7_io_outputC[25:0]     ), //o
    .clk                     (clk                          ), //i
    .reset                   (reset                        )  //i
  );
  ProcessingElement pes_0_8 (
    .io_inputA               (pes_0_7_io_outputA[7:0]      ), //i
    .io_inputB               (skewBuffer_1_io_output_8[7:0]), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_0_8  ), //i
    .io_resetPartialC        (io_resetPartialC_0_8         ), //i
    .io_outputA              (pes_0_8_io_outputA[7:0]      ), //o
    .io_outputB              (pes_0_8_io_outputB[7:0]      ), //o
    .io_outputC              (pes_0_8_io_outputC[25:0]     ), //o
    .clk                     (clk                          ), //i
    .reset                   (reset                        )  //i
  );
  ProcessingElement pes_0_9 (
    .io_inputA               (pes_0_8_io_outputA[7:0]      ), //i
    .io_inputB               (skewBuffer_1_io_output_9[7:0]), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_0_9  ), //i
    .io_resetPartialC        (io_resetPartialC_0_9         ), //i
    .io_outputA              (pes_0_9_io_outputA[7:0]      ), //o
    .io_outputB              (pes_0_9_io_outputB[7:0]      ), //o
    .io_outputC              (pes_0_9_io_outputC[25:0]     ), //o
    .clk                     (clk                          ), //i
    .reset                   (reset                        )  //i
  );
  ProcessingElement pes_0_10 (
    .io_inputA               (pes_0_9_io_outputA[7:0]       ), //i
    .io_inputB               (skewBuffer_1_io_output_10[7:0]), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_0_10  ), //i
    .io_resetPartialC        (io_resetPartialC_0_10         ), //i
    .io_outputA              (pes_0_10_io_outputA[7:0]      ), //o
    .io_outputB              (pes_0_10_io_outputB[7:0]      ), //o
    .io_outputC              (pes_0_10_io_outputC[25:0]     ), //o
    .clk                     (clk                           ), //i
    .reset                   (reset                         )  //i
  );
  ProcessingElement pes_0_11 (
    .io_inputA               (pes_0_10_io_outputA[7:0]      ), //i
    .io_inputB               (skewBuffer_1_io_output_11[7:0]), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_0_11  ), //i
    .io_resetPartialC        (io_resetPartialC_0_11         ), //i
    .io_outputA              (pes_0_11_io_outputA[7:0]      ), //o
    .io_outputB              (pes_0_11_io_outputB[7:0]      ), //o
    .io_outputC              (pes_0_11_io_outputC[25:0]     ), //o
    .clk                     (clk                           ), //i
    .reset                   (reset                         )  //i
  );
  ProcessingElement pes_0_12 (
    .io_inputA               (pes_0_11_io_outputA[7:0]      ), //i
    .io_inputB               (skewBuffer_1_io_output_12[7:0]), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_0_12  ), //i
    .io_resetPartialC        (io_resetPartialC_0_12         ), //i
    .io_outputA              (pes_0_12_io_outputA[7:0]      ), //o
    .io_outputB              (pes_0_12_io_outputB[7:0]      ), //o
    .io_outputC              (pes_0_12_io_outputC[25:0]     ), //o
    .clk                     (clk                           ), //i
    .reset                   (reset                         )  //i
  );
  ProcessingElement pes_0_13 (
    .io_inputA               (pes_0_12_io_outputA[7:0]      ), //i
    .io_inputB               (skewBuffer_1_io_output_13[7:0]), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_0_13  ), //i
    .io_resetPartialC        (io_resetPartialC_0_13         ), //i
    .io_outputA              (pes_0_13_io_outputA[7:0]      ), //o
    .io_outputB              (pes_0_13_io_outputB[7:0]      ), //o
    .io_outputC              (pes_0_13_io_outputC[25:0]     ), //o
    .clk                     (clk                           ), //i
    .reset                   (reset                         )  //i
  );
  ProcessingElement pes_0_14 (
    .io_inputA               (pes_0_13_io_outputA[7:0]      ), //i
    .io_inputB               (skewBuffer_1_io_output_14[7:0]), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_0_14  ), //i
    .io_resetPartialC        (io_resetPartialC_0_14         ), //i
    .io_outputA              (pes_0_14_io_outputA[7:0]      ), //o
    .io_outputB              (pes_0_14_io_outputB[7:0]      ), //o
    .io_outputC              (pes_0_14_io_outputC[25:0]     ), //o
    .clk                     (clk                           ), //i
    .reset                   (reset                         )  //i
  );
  ProcessingElement_15 pes_0_15 (
    .io_inputA               (pes_0_14_io_outputA[7:0]      ), //i
    .io_inputB               (skewBuffer_1_io_output_15[7:0]), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_0_15  ), //i
    .io_resetPartialC        (io_resetPartialC_0_15         ), //i
    .io_outputB              (pes_0_15_io_outputB[7:0]      ), //o
    .io_outputC              (pes_0_15_io_outputC[25:0]     ), //o
    .clk                     (clk                           ), //i
    .reset                   (reset                         )  //i
  );
  ProcessingElement_16 pes_1_0 (
    .io_inputA               (skewBuffer_io_output_1[7:0]), //i
    .io_inputB               (pes_0_0_io_outputB[7:0]    ), //i
    .io_inputC               (pes_0_1_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_1_0), //i
    .io_resetPartialC        (io_resetPartialC_1_0       ), //i
    .io_outputA              (pes_1_0_io_outputA[7:0]    ), //o
    .io_outputB              (pes_1_0_io_outputB[7:0]    ), //o
    .io_outputC              (pes_1_0_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_1_1 (
    .io_inputA               (pes_1_0_io_outputA[7:0]    ), //i
    .io_inputB               (pes_0_1_io_outputB[7:0]    ), //i
    .io_inputC               (pes_0_2_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_1_1), //i
    .io_resetPartialC        (io_resetPartialC_1_1       ), //i
    .io_outputA              (pes_1_1_io_outputA[7:0]    ), //o
    .io_outputB              (pes_1_1_io_outputB[7:0]    ), //o
    .io_outputC              (pes_1_1_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_1_2 (
    .io_inputA               (pes_1_1_io_outputA[7:0]    ), //i
    .io_inputB               (pes_0_2_io_outputB[7:0]    ), //i
    .io_inputC               (pes_0_3_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_1_2), //i
    .io_resetPartialC        (io_resetPartialC_1_2       ), //i
    .io_outputA              (pes_1_2_io_outputA[7:0]    ), //o
    .io_outputB              (pes_1_2_io_outputB[7:0]    ), //o
    .io_outputC              (pes_1_2_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_1_3 (
    .io_inputA               (pes_1_2_io_outputA[7:0]    ), //i
    .io_inputB               (pes_0_3_io_outputB[7:0]    ), //i
    .io_inputC               (pes_0_4_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_1_3), //i
    .io_resetPartialC        (io_resetPartialC_1_3       ), //i
    .io_outputA              (pes_1_3_io_outputA[7:0]    ), //o
    .io_outputB              (pes_1_3_io_outputB[7:0]    ), //o
    .io_outputC              (pes_1_3_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_1_4 (
    .io_inputA               (pes_1_3_io_outputA[7:0]    ), //i
    .io_inputB               (pes_0_4_io_outputB[7:0]    ), //i
    .io_inputC               (pes_0_5_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_1_4), //i
    .io_resetPartialC        (io_resetPartialC_1_4       ), //i
    .io_outputA              (pes_1_4_io_outputA[7:0]    ), //o
    .io_outputB              (pes_1_4_io_outputB[7:0]    ), //o
    .io_outputC              (pes_1_4_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_1_5 (
    .io_inputA               (pes_1_4_io_outputA[7:0]    ), //i
    .io_inputB               (pes_0_5_io_outputB[7:0]    ), //i
    .io_inputC               (pes_0_6_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_1_5), //i
    .io_resetPartialC        (io_resetPartialC_1_5       ), //i
    .io_outputA              (pes_1_5_io_outputA[7:0]    ), //o
    .io_outputB              (pes_1_5_io_outputB[7:0]    ), //o
    .io_outputC              (pes_1_5_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_1_6 (
    .io_inputA               (pes_1_5_io_outputA[7:0]    ), //i
    .io_inputB               (pes_0_6_io_outputB[7:0]    ), //i
    .io_inputC               (pes_0_7_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_1_6), //i
    .io_resetPartialC        (io_resetPartialC_1_6       ), //i
    .io_outputA              (pes_1_6_io_outputA[7:0]    ), //o
    .io_outputB              (pes_1_6_io_outputB[7:0]    ), //o
    .io_outputC              (pes_1_6_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_1_7 (
    .io_inputA               (pes_1_6_io_outputA[7:0]    ), //i
    .io_inputB               (pes_0_7_io_outputB[7:0]    ), //i
    .io_inputC               (pes_0_8_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_1_7), //i
    .io_resetPartialC        (io_resetPartialC_1_7       ), //i
    .io_outputA              (pes_1_7_io_outputA[7:0]    ), //o
    .io_outputB              (pes_1_7_io_outputB[7:0]    ), //o
    .io_outputC              (pes_1_7_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_1_8 (
    .io_inputA               (pes_1_7_io_outputA[7:0]    ), //i
    .io_inputB               (pes_0_8_io_outputB[7:0]    ), //i
    .io_inputC               (pes_0_9_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_1_8), //i
    .io_resetPartialC        (io_resetPartialC_1_8       ), //i
    .io_outputA              (pes_1_8_io_outputA[7:0]    ), //o
    .io_outputB              (pes_1_8_io_outputB[7:0]    ), //o
    .io_outputC              (pes_1_8_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_1_9 (
    .io_inputA               (pes_1_8_io_outputA[7:0]    ), //i
    .io_inputB               (pes_0_9_io_outputB[7:0]    ), //i
    .io_inputC               (pes_0_10_io_outputC[25:0]  ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_1_9), //i
    .io_resetPartialC        (io_resetPartialC_1_9       ), //i
    .io_outputA              (pes_1_9_io_outputA[7:0]    ), //o
    .io_outputB              (pes_1_9_io_outputB[7:0]    ), //o
    .io_outputC              (pes_1_9_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_1_10 (
    .io_inputA               (pes_1_9_io_outputA[7:0]     ), //i
    .io_inputB               (pes_0_10_io_outputB[7:0]    ), //i
    .io_inputC               (pes_0_11_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_1_10), //i
    .io_resetPartialC        (io_resetPartialC_1_10       ), //i
    .io_outputA              (pes_1_10_io_outputA[7:0]    ), //o
    .io_outputB              (pes_1_10_io_outputB[7:0]    ), //o
    .io_outputC              (pes_1_10_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_1_11 (
    .io_inputA               (pes_1_10_io_outputA[7:0]    ), //i
    .io_inputB               (pes_0_11_io_outputB[7:0]    ), //i
    .io_inputC               (pes_0_12_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_1_11), //i
    .io_resetPartialC        (io_resetPartialC_1_11       ), //i
    .io_outputA              (pes_1_11_io_outputA[7:0]    ), //o
    .io_outputB              (pes_1_11_io_outputB[7:0]    ), //o
    .io_outputC              (pes_1_11_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_1_12 (
    .io_inputA               (pes_1_11_io_outputA[7:0]    ), //i
    .io_inputB               (pes_0_12_io_outputB[7:0]    ), //i
    .io_inputC               (pes_0_13_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_1_12), //i
    .io_resetPartialC        (io_resetPartialC_1_12       ), //i
    .io_outputA              (pes_1_12_io_outputA[7:0]    ), //o
    .io_outputB              (pes_1_12_io_outputB[7:0]    ), //o
    .io_outputC              (pes_1_12_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_1_13 (
    .io_inputA               (pes_1_12_io_outputA[7:0]    ), //i
    .io_inputB               (pes_0_13_io_outputB[7:0]    ), //i
    .io_inputC               (pes_0_14_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_1_13), //i
    .io_resetPartialC        (io_resetPartialC_1_13       ), //i
    .io_outputA              (pes_1_13_io_outputA[7:0]    ), //o
    .io_outputB              (pes_1_13_io_outputB[7:0]    ), //o
    .io_outputC              (pes_1_13_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_1_14 (
    .io_inputA               (pes_1_13_io_outputA[7:0]    ), //i
    .io_inputB               (pes_0_14_io_outputB[7:0]    ), //i
    .io_inputC               (pes_0_15_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_1_14), //i
    .io_resetPartialC        (io_resetPartialC_1_14       ), //i
    .io_outputA              (pes_1_14_io_outputA[7:0]    ), //o
    .io_outputB              (pes_1_14_io_outputB[7:0]    ), //o
    .io_outputC              (pes_1_14_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_15 pes_1_15 (
    .io_inputA               (pes_1_14_io_outputA[7:0]    ), //i
    .io_inputB               (pes_0_15_io_outputB[7:0]    ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_1_15), //i
    .io_resetPartialC        (io_resetPartialC_1_15       ), //i
    .io_outputB              (pes_1_15_io_outputB[7:0]    ), //o
    .io_outputC              (pes_1_15_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_2_0 (
    .io_inputA               (skewBuffer_io_output_2[7:0]), //i
    .io_inputB               (pes_1_0_io_outputB[7:0]    ), //i
    .io_inputC               (pes_1_1_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_2_0), //i
    .io_resetPartialC        (io_resetPartialC_2_0       ), //i
    .io_outputA              (pes_2_0_io_outputA[7:0]    ), //o
    .io_outputB              (pes_2_0_io_outputB[7:0]    ), //o
    .io_outputC              (pes_2_0_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_2_1 (
    .io_inputA               (pes_2_0_io_outputA[7:0]    ), //i
    .io_inputB               (pes_1_1_io_outputB[7:0]    ), //i
    .io_inputC               (pes_1_2_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_2_1), //i
    .io_resetPartialC        (io_resetPartialC_2_1       ), //i
    .io_outputA              (pes_2_1_io_outputA[7:0]    ), //o
    .io_outputB              (pes_2_1_io_outputB[7:0]    ), //o
    .io_outputC              (pes_2_1_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_2_2 (
    .io_inputA               (pes_2_1_io_outputA[7:0]    ), //i
    .io_inputB               (pes_1_2_io_outputB[7:0]    ), //i
    .io_inputC               (pes_1_3_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_2_2), //i
    .io_resetPartialC        (io_resetPartialC_2_2       ), //i
    .io_outputA              (pes_2_2_io_outputA[7:0]    ), //o
    .io_outputB              (pes_2_2_io_outputB[7:0]    ), //o
    .io_outputC              (pes_2_2_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_2_3 (
    .io_inputA               (pes_2_2_io_outputA[7:0]    ), //i
    .io_inputB               (pes_1_3_io_outputB[7:0]    ), //i
    .io_inputC               (pes_1_4_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_2_3), //i
    .io_resetPartialC        (io_resetPartialC_2_3       ), //i
    .io_outputA              (pes_2_3_io_outputA[7:0]    ), //o
    .io_outputB              (pes_2_3_io_outputB[7:0]    ), //o
    .io_outputC              (pes_2_3_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_2_4 (
    .io_inputA               (pes_2_3_io_outputA[7:0]    ), //i
    .io_inputB               (pes_1_4_io_outputB[7:0]    ), //i
    .io_inputC               (pes_1_5_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_2_4), //i
    .io_resetPartialC        (io_resetPartialC_2_4       ), //i
    .io_outputA              (pes_2_4_io_outputA[7:0]    ), //o
    .io_outputB              (pes_2_4_io_outputB[7:0]    ), //o
    .io_outputC              (pes_2_4_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_2_5 (
    .io_inputA               (pes_2_4_io_outputA[7:0]    ), //i
    .io_inputB               (pes_1_5_io_outputB[7:0]    ), //i
    .io_inputC               (pes_1_6_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_2_5), //i
    .io_resetPartialC        (io_resetPartialC_2_5       ), //i
    .io_outputA              (pes_2_5_io_outputA[7:0]    ), //o
    .io_outputB              (pes_2_5_io_outputB[7:0]    ), //o
    .io_outputC              (pes_2_5_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_2_6 (
    .io_inputA               (pes_2_5_io_outputA[7:0]    ), //i
    .io_inputB               (pes_1_6_io_outputB[7:0]    ), //i
    .io_inputC               (pes_1_7_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_2_6), //i
    .io_resetPartialC        (io_resetPartialC_2_6       ), //i
    .io_outputA              (pes_2_6_io_outputA[7:0]    ), //o
    .io_outputB              (pes_2_6_io_outputB[7:0]    ), //o
    .io_outputC              (pes_2_6_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_2_7 (
    .io_inputA               (pes_2_6_io_outputA[7:0]    ), //i
    .io_inputB               (pes_1_7_io_outputB[7:0]    ), //i
    .io_inputC               (pes_1_8_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_2_7), //i
    .io_resetPartialC        (io_resetPartialC_2_7       ), //i
    .io_outputA              (pes_2_7_io_outputA[7:0]    ), //o
    .io_outputB              (pes_2_7_io_outputB[7:0]    ), //o
    .io_outputC              (pes_2_7_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_2_8 (
    .io_inputA               (pes_2_7_io_outputA[7:0]    ), //i
    .io_inputB               (pes_1_8_io_outputB[7:0]    ), //i
    .io_inputC               (pes_1_9_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_2_8), //i
    .io_resetPartialC        (io_resetPartialC_2_8       ), //i
    .io_outputA              (pes_2_8_io_outputA[7:0]    ), //o
    .io_outputB              (pes_2_8_io_outputB[7:0]    ), //o
    .io_outputC              (pes_2_8_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_2_9 (
    .io_inputA               (pes_2_8_io_outputA[7:0]    ), //i
    .io_inputB               (pes_1_9_io_outputB[7:0]    ), //i
    .io_inputC               (pes_1_10_io_outputC[25:0]  ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_2_9), //i
    .io_resetPartialC        (io_resetPartialC_2_9       ), //i
    .io_outputA              (pes_2_9_io_outputA[7:0]    ), //o
    .io_outputB              (pes_2_9_io_outputB[7:0]    ), //o
    .io_outputC              (pes_2_9_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_2_10 (
    .io_inputA               (pes_2_9_io_outputA[7:0]     ), //i
    .io_inputB               (pes_1_10_io_outputB[7:0]    ), //i
    .io_inputC               (pes_1_11_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_2_10), //i
    .io_resetPartialC        (io_resetPartialC_2_10       ), //i
    .io_outputA              (pes_2_10_io_outputA[7:0]    ), //o
    .io_outputB              (pes_2_10_io_outputB[7:0]    ), //o
    .io_outputC              (pes_2_10_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_2_11 (
    .io_inputA               (pes_2_10_io_outputA[7:0]    ), //i
    .io_inputB               (pes_1_11_io_outputB[7:0]    ), //i
    .io_inputC               (pes_1_12_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_2_11), //i
    .io_resetPartialC        (io_resetPartialC_2_11       ), //i
    .io_outputA              (pes_2_11_io_outputA[7:0]    ), //o
    .io_outputB              (pes_2_11_io_outputB[7:0]    ), //o
    .io_outputC              (pes_2_11_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_2_12 (
    .io_inputA               (pes_2_11_io_outputA[7:0]    ), //i
    .io_inputB               (pes_1_12_io_outputB[7:0]    ), //i
    .io_inputC               (pes_1_13_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_2_12), //i
    .io_resetPartialC        (io_resetPartialC_2_12       ), //i
    .io_outputA              (pes_2_12_io_outputA[7:0]    ), //o
    .io_outputB              (pes_2_12_io_outputB[7:0]    ), //o
    .io_outputC              (pes_2_12_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_2_13 (
    .io_inputA               (pes_2_12_io_outputA[7:0]    ), //i
    .io_inputB               (pes_1_13_io_outputB[7:0]    ), //i
    .io_inputC               (pes_1_14_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_2_13), //i
    .io_resetPartialC        (io_resetPartialC_2_13       ), //i
    .io_outputA              (pes_2_13_io_outputA[7:0]    ), //o
    .io_outputB              (pes_2_13_io_outputB[7:0]    ), //o
    .io_outputC              (pes_2_13_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_2_14 (
    .io_inputA               (pes_2_13_io_outputA[7:0]    ), //i
    .io_inputB               (pes_1_14_io_outputB[7:0]    ), //i
    .io_inputC               (pes_1_15_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_2_14), //i
    .io_resetPartialC        (io_resetPartialC_2_14       ), //i
    .io_outputA              (pes_2_14_io_outputA[7:0]    ), //o
    .io_outputB              (pes_2_14_io_outputB[7:0]    ), //o
    .io_outputC              (pes_2_14_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_15 pes_2_15 (
    .io_inputA               (pes_2_14_io_outputA[7:0]    ), //i
    .io_inputB               (pes_1_15_io_outputB[7:0]    ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_2_15), //i
    .io_resetPartialC        (io_resetPartialC_2_15       ), //i
    .io_outputB              (pes_2_15_io_outputB[7:0]    ), //o
    .io_outputC              (pes_2_15_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_3_0 (
    .io_inputA               (skewBuffer_io_output_3[7:0]), //i
    .io_inputB               (pes_2_0_io_outputB[7:0]    ), //i
    .io_inputC               (pes_2_1_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_3_0), //i
    .io_resetPartialC        (io_resetPartialC_3_0       ), //i
    .io_outputA              (pes_3_0_io_outputA[7:0]    ), //o
    .io_outputB              (pes_3_0_io_outputB[7:0]    ), //o
    .io_outputC              (pes_3_0_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_3_1 (
    .io_inputA               (pes_3_0_io_outputA[7:0]    ), //i
    .io_inputB               (pes_2_1_io_outputB[7:0]    ), //i
    .io_inputC               (pes_2_2_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_3_1), //i
    .io_resetPartialC        (io_resetPartialC_3_1       ), //i
    .io_outputA              (pes_3_1_io_outputA[7:0]    ), //o
    .io_outputB              (pes_3_1_io_outputB[7:0]    ), //o
    .io_outputC              (pes_3_1_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_3_2 (
    .io_inputA               (pes_3_1_io_outputA[7:0]    ), //i
    .io_inputB               (pes_2_2_io_outputB[7:0]    ), //i
    .io_inputC               (pes_2_3_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_3_2), //i
    .io_resetPartialC        (io_resetPartialC_3_2       ), //i
    .io_outputA              (pes_3_2_io_outputA[7:0]    ), //o
    .io_outputB              (pes_3_2_io_outputB[7:0]    ), //o
    .io_outputC              (pes_3_2_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_3_3 (
    .io_inputA               (pes_3_2_io_outputA[7:0]    ), //i
    .io_inputB               (pes_2_3_io_outputB[7:0]    ), //i
    .io_inputC               (pes_2_4_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_3_3), //i
    .io_resetPartialC        (io_resetPartialC_3_3       ), //i
    .io_outputA              (pes_3_3_io_outputA[7:0]    ), //o
    .io_outputB              (pes_3_3_io_outputB[7:0]    ), //o
    .io_outputC              (pes_3_3_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_3_4 (
    .io_inputA               (pes_3_3_io_outputA[7:0]    ), //i
    .io_inputB               (pes_2_4_io_outputB[7:0]    ), //i
    .io_inputC               (pes_2_5_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_3_4), //i
    .io_resetPartialC        (io_resetPartialC_3_4       ), //i
    .io_outputA              (pes_3_4_io_outputA[7:0]    ), //o
    .io_outputB              (pes_3_4_io_outputB[7:0]    ), //o
    .io_outputC              (pes_3_4_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_3_5 (
    .io_inputA               (pes_3_4_io_outputA[7:0]    ), //i
    .io_inputB               (pes_2_5_io_outputB[7:0]    ), //i
    .io_inputC               (pes_2_6_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_3_5), //i
    .io_resetPartialC        (io_resetPartialC_3_5       ), //i
    .io_outputA              (pes_3_5_io_outputA[7:0]    ), //o
    .io_outputB              (pes_3_5_io_outputB[7:0]    ), //o
    .io_outputC              (pes_3_5_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_3_6 (
    .io_inputA               (pes_3_5_io_outputA[7:0]    ), //i
    .io_inputB               (pes_2_6_io_outputB[7:0]    ), //i
    .io_inputC               (pes_2_7_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_3_6), //i
    .io_resetPartialC        (io_resetPartialC_3_6       ), //i
    .io_outputA              (pes_3_6_io_outputA[7:0]    ), //o
    .io_outputB              (pes_3_6_io_outputB[7:0]    ), //o
    .io_outputC              (pes_3_6_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_3_7 (
    .io_inputA               (pes_3_6_io_outputA[7:0]    ), //i
    .io_inputB               (pes_2_7_io_outputB[7:0]    ), //i
    .io_inputC               (pes_2_8_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_3_7), //i
    .io_resetPartialC        (io_resetPartialC_3_7       ), //i
    .io_outputA              (pes_3_7_io_outputA[7:0]    ), //o
    .io_outputB              (pes_3_7_io_outputB[7:0]    ), //o
    .io_outputC              (pes_3_7_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_3_8 (
    .io_inputA               (pes_3_7_io_outputA[7:0]    ), //i
    .io_inputB               (pes_2_8_io_outputB[7:0]    ), //i
    .io_inputC               (pes_2_9_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_3_8), //i
    .io_resetPartialC        (io_resetPartialC_3_8       ), //i
    .io_outputA              (pes_3_8_io_outputA[7:0]    ), //o
    .io_outputB              (pes_3_8_io_outputB[7:0]    ), //o
    .io_outputC              (pes_3_8_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_3_9 (
    .io_inputA               (pes_3_8_io_outputA[7:0]    ), //i
    .io_inputB               (pes_2_9_io_outputB[7:0]    ), //i
    .io_inputC               (pes_2_10_io_outputC[25:0]  ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_3_9), //i
    .io_resetPartialC        (io_resetPartialC_3_9       ), //i
    .io_outputA              (pes_3_9_io_outputA[7:0]    ), //o
    .io_outputB              (pes_3_9_io_outputB[7:0]    ), //o
    .io_outputC              (pes_3_9_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_3_10 (
    .io_inputA               (pes_3_9_io_outputA[7:0]     ), //i
    .io_inputB               (pes_2_10_io_outputB[7:0]    ), //i
    .io_inputC               (pes_2_11_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_3_10), //i
    .io_resetPartialC        (io_resetPartialC_3_10       ), //i
    .io_outputA              (pes_3_10_io_outputA[7:0]    ), //o
    .io_outputB              (pes_3_10_io_outputB[7:0]    ), //o
    .io_outputC              (pes_3_10_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_3_11 (
    .io_inputA               (pes_3_10_io_outputA[7:0]    ), //i
    .io_inputB               (pes_2_11_io_outputB[7:0]    ), //i
    .io_inputC               (pes_2_12_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_3_11), //i
    .io_resetPartialC        (io_resetPartialC_3_11       ), //i
    .io_outputA              (pes_3_11_io_outputA[7:0]    ), //o
    .io_outputB              (pes_3_11_io_outputB[7:0]    ), //o
    .io_outputC              (pes_3_11_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_3_12 (
    .io_inputA               (pes_3_11_io_outputA[7:0]    ), //i
    .io_inputB               (pes_2_12_io_outputB[7:0]    ), //i
    .io_inputC               (pes_2_13_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_3_12), //i
    .io_resetPartialC        (io_resetPartialC_3_12       ), //i
    .io_outputA              (pes_3_12_io_outputA[7:0]    ), //o
    .io_outputB              (pes_3_12_io_outputB[7:0]    ), //o
    .io_outputC              (pes_3_12_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_3_13 (
    .io_inputA               (pes_3_12_io_outputA[7:0]    ), //i
    .io_inputB               (pes_2_13_io_outputB[7:0]    ), //i
    .io_inputC               (pes_2_14_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_3_13), //i
    .io_resetPartialC        (io_resetPartialC_3_13       ), //i
    .io_outputA              (pes_3_13_io_outputA[7:0]    ), //o
    .io_outputB              (pes_3_13_io_outputB[7:0]    ), //o
    .io_outputC              (pes_3_13_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_3_14 (
    .io_inputA               (pes_3_13_io_outputA[7:0]    ), //i
    .io_inputB               (pes_2_14_io_outputB[7:0]    ), //i
    .io_inputC               (pes_2_15_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_3_14), //i
    .io_resetPartialC        (io_resetPartialC_3_14       ), //i
    .io_outputA              (pes_3_14_io_outputA[7:0]    ), //o
    .io_outputB              (pes_3_14_io_outputB[7:0]    ), //o
    .io_outputC              (pes_3_14_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_15 pes_3_15 (
    .io_inputA               (pes_3_14_io_outputA[7:0]    ), //i
    .io_inputB               (pes_2_15_io_outputB[7:0]    ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_3_15), //i
    .io_resetPartialC        (io_resetPartialC_3_15       ), //i
    .io_outputB              (pes_3_15_io_outputB[7:0]    ), //o
    .io_outputC              (pes_3_15_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_4_0 (
    .io_inputA               (skewBuffer_io_output_4[7:0]), //i
    .io_inputB               (pes_3_0_io_outputB[7:0]    ), //i
    .io_inputC               (pes_3_1_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_4_0), //i
    .io_resetPartialC        (io_resetPartialC_4_0       ), //i
    .io_outputA              (pes_4_0_io_outputA[7:0]    ), //o
    .io_outputB              (pes_4_0_io_outputB[7:0]    ), //o
    .io_outputC              (pes_4_0_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_4_1 (
    .io_inputA               (pes_4_0_io_outputA[7:0]    ), //i
    .io_inputB               (pes_3_1_io_outputB[7:0]    ), //i
    .io_inputC               (pes_3_2_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_4_1), //i
    .io_resetPartialC        (io_resetPartialC_4_1       ), //i
    .io_outputA              (pes_4_1_io_outputA[7:0]    ), //o
    .io_outputB              (pes_4_1_io_outputB[7:0]    ), //o
    .io_outputC              (pes_4_1_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_4_2 (
    .io_inputA               (pes_4_1_io_outputA[7:0]    ), //i
    .io_inputB               (pes_3_2_io_outputB[7:0]    ), //i
    .io_inputC               (pes_3_3_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_4_2), //i
    .io_resetPartialC        (io_resetPartialC_4_2       ), //i
    .io_outputA              (pes_4_2_io_outputA[7:0]    ), //o
    .io_outputB              (pes_4_2_io_outputB[7:0]    ), //o
    .io_outputC              (pes_4_2_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_4_3 (
    .io_inputA               (pes_4_2_io_outputA[7:0]    ), //i
    .io_inputB               (pes_3_3_io_outputB[7:0]    ), //i
    .io_inputC               (pes_3_4_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_4_3), //i
    .io_resetPartialC        (io_resetPartialC_4_3       ), //i
    .io_outputA              (pes_4_3_io_outputA[7:0]    ), //o
    .io_outputB              (pes_4_3_io_outputB[7:0]    ), //o
    .io_outputC              (pes_4_3_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_4_4 (
    .io_inputA               (pes_4_3_io_outputA[7:0]    ), //i
    .io_inputB               (pes_3_4_io_outputB[7:0]    ), //i
    .io_inputC               (pes_3_5_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_4_4), //i
    .io_resetPartialC        (io_resetPartialC_4_4       ), //i
    .io_outputA              (pes_4_4_io_outputA[7:0]    ), //o
    .io_outputB              (pes_4_4_io_outputB[7:0]    ), //o
    .io_outputC              (pes_4_4_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_4_5 (
    .io_inputA               (pes_4_4_io_outputA[7:0]    ), //i
    .io_inputB               (pes_3_5_io_outputB[7:0]    ), //i
    .io_inputC               (pes_3_6_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_4_5), //i
    .io_resetPartialC        (io_resetPartialC_4_5       ), //i
    .io_outputA              (pes_4_5_io_outputA[7:0]    ), //o
    .io_outputB              (pes_4_5_io_outputB[7:0]    ), //o
    .io_outputC              (pes_4_5_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_4_6 (
    .io_inputA               (pes_4_5_io_outputA[7:0]    ), //i
    .io_inputB               (pes_3_6_io_outputB[7:0]    ), //i
    .io_inputC               (pes_3_7_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_4_6), //i
    .io_resetPartialC        (io_resetPartialC_4_6       ), //i
    .io_outputA              (pes_4_6_io_outputA[7:0]    ), //o
    .io_outputB              (pes_4_6_io_outputB[7:0]    ), //o
    .io_outputC              (pes_4_6_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_4_7 (
    .io_inputA               (pes_4_6_io_outputA[7:0]    ), //i
    .io_inputB               (pes_3_7_io_outputB[7:0]    ), //i
    .io_inputC               (pes_3_8_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_4_7), //i
    .io_resetPartialC        (io_resetPartialC_4_7       ), //i
    .io_outputA              (pes_4_7_io_outputA[7:0]    ), //o
    .io_outputB              (pes_4_7_io_outputB[7:0]    ), //o
    .io_outputC              (pes_4_7_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_4_8 (
    .io_inputA               (pes_4_7_io_outputA[7:0]    ), //i
    .io_inputB               (pes_3_8_io_outputB[7:0]    ), //i
    .io_inputC               (pes_3_9_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_4_8), //i
    .io_resetPartialC        (io_resetPartialC_4_8       ), //i
    .io_outputA              (pes_4_8_io_outputA[7:0]    ), //o
    .io_outputB              (pes_4_8_io_outputB[7:0]    ), //o
    .io_outputC              (pes_4_8_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_4_9 (
    .io_inputA               (pes_4_8_io_outputA[7:0]    ), //i
    .io_inputB               (pes_3_9_io_outputB[7:0]    ), //i
    .io_inputC               (pes_3_10_io_outputC[25:0]  ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_4_9), //i
    .io_resetPartialC        (io_resetPartialC_4_9       ), //i
    .io_outputA              (pes_4_9_io_outputA[7:0]    ), //o
    .io_outputB              (pes_4_9_io_outputB[7:0]    ), //o
    .io_outputC              (pes_4_9_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_4_10 (
    .io_inputA               (pes_4_9_io_outputA[7:0]     ), //i
    .io_inputB               (pes_3_10_io_outputB[7:0]    ), //i
    .io_inputC               (pes_3_11_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_4_10), //i
    .io_resetPartialC        (io_resetPartialC_4_10       ), //i
    .io_outputA              (pes_4_10_io_outputA[7:0]    ), //o
    .io_outputB              (pes_4_10_io_outputB[7:0]    ), //o
    .io_outputC              (pes_4_10_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_4_11 (
    .io_inputA               (pes_4_10_io_outputA[7:0]    ), //i
    .io_inputB               (pes_3_11_io_outputB[7:0]    ), //i
    .io_inputC               (pes_3_12_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_4_11), //i
    .io_resetPartialC        (io_resetPartialC_4_11       ), //i
    .io_outputA              (pes_4_11_io_outputA[7:0]    ), //o
    .io_outputB              (pes_4_11_io_outputB[7:0]    ), //o
    .io_outputC              (pes_4_11_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_4_12 (
    .io_inputA               (pes_4_11_io_outputA[7:0]    ), //i
    .io_inputB               (pes_3_12_io_outputB[7:0]    ), //i
    .io_inputC               (pes_3_13_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_4_12), //i
    .io_resetPartialC        (io_resetPartialC_4_12       ), //i
    .io_outputA              (pes_4_12_io_outputA[7:0]    ), //o
    .io_outputB              (pes_4_12_io_outputB[7:0]    ), //o
    .io_outputC              (pes_4_12_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_4_13 (
    .io_inputA               (pes_4_12_io_outputA[7:0]    ), //i
    .io_inputB               (pes_3_13_io_outputB[7:0]    ), //i
    .io_inputC               (pes_3_14_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_4_13), //i
    .io_resetPartialC        (io_resetPartialC_4_13       ), //i
    .io_outputA              (pes_4_13_io_outputA[7:0]    ), //o
    .io_outputB              (pes_4_13_io_outputB[7:0]    ), //o
    .io_outputC              (pes_4_13_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_4_14 (
    .io_inputA               (pes_4_13_io_outputA[7:0]    ), //i
    .io_inputB               (pes_3_14_io_outputB[7:0]    ), //i
    .io_inputC               (pes_3_15_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_4_14), //i
    .io_resetPartialC        (io_resetPartialC_4_14       ), //i
    .io_outputA              (pes_4_14_io_outputA[7:0]    ), //o
    .io_outputB              (pes_4_14_io_outputB[7:0]    ), //o
    .io_outputC              (pes_4_14_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_15 pes_4_15 (
    .io_inputA               (pes_4_14_io_outputA[7:0]    ), //i
    .io_inputB               (pes_3_15_io_outputB[7:0]    ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_4_15), //i
    .io_resetPartialC        (io_resetPartialC_4_15       ), //i
    .io_outputB              (pes_4_15_io_outputB[7:0]    ), //o
    .io_outputC              (pes_4_15_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_5_0 (
    .io_inputA               (skewBuffer_io_output_5[7:0]), //i
    .io_inputB               (pes_4_0_io_outputB[7:0]    ), //i
    .io_inputC               (pes_4_1_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_5_0), //i
    .io_resetPartialC        (io_resetPartialC_5_0       ), //i
    .io_outputA              (pes_5_0_io_outputA[7:0]    ), //o
    .io_outputB              (pes_5_0_io_outputB[7:0]    ), //o
    .io_outputC              (pes_5_0_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_5_1 (
    .io_inputA               (pes_5_0_io_outputA[7:0]    ), //i
    .io_inputB               (pes_4_1_io_outputB[7:0]    ), //i
    .io_inputC               (pes_4_2_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_5_1), //i
    .io_resetPartialC        (io_resetPartialC_5_1       ), //i
    .io_outputA              (pes_5_1_io_outputA[7:0]    ), //o
    .io_outputB              (pes_5_1_io_outputB[7:0]    ), //o
    .io_outputC              (pes_5_1_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_5_2 (
    .io_inputA               (pes_5_1_io_outputA[7:0]    ), //i
    .io_inputB               (pes_4_2_io_outputB[7:0]    ), //i
    .io_inputC               (pes_4_3_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_5_2), //i
    .io_resetPartialC        (io_resetPartialC_5_2       ), //i
    .io_outputA              (pes_5_2_io_outputA[7:0]    ), //o
    .io_outputB              (pes_5_2_io_outputB[7:0]    ), //o
    .io_outputC              (pes_5_2_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_5_3 (
    .io_inputA               (pes_5_2_io_outputA[7:0]    ), //i
    .io_inputB               (pes_4_3_io_outputB[7:0]    ), //i
    .io_inputC               (pes_4_4_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_5_3), //i
    .io_resetPartialC        (io_resetPartialC_5_3       ), //i
    .io_outputA              (pes_5_3_io_outputA[7:0]    ), //o
    .io_outputB              (pes_5_3_io_outputB[7:0]    ), //o
    .io_outputC              (pes_5_3_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_5_4 (
    .io_inputA               (pes_5_3_io_outputA[7:0]    ), //i
    .io_inputB               (pes_4_4_io_outputB[7:0]    ), //i
    .io_inputC               (pes_4_5_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_5_4), //i
    .io_resetPartialC        (io_resetPartialC_5_4       ), //i
    .io_outputA              (pes_5_4_io_outputA[7:0]    ), //o
    .io_outputB              (pes_5_4_io_outputB[7:0]    ), //o
    .io_outputC              (pes_5_4_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_5_5 (
    .io_inputA               (pes_5_4_io_outputA[7:0]    ), //i
    .io_inputB               (pes_4_5_io_outputB[7:0]    ), //i
    .io_inputC               (pes_4_6_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_5_5), //i
    .io_resetPartialC        (io_resetPartialC_5_5       ), //i
    .io_outputA              (pes_5_5_io_outputA[7:0]    ), //o
    .io_outputB              (pes_5_5_io_outputB[7:0]    ), //o
    .io_outputC              (pes_5_5_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_5_6 (
    .io_inputA               (pes_5_5_io_outputA[7:0]    ), //i
    .io_inputB               (pes_4_6_io_outputB[7:0]    ), //i
    .io_inputC               (pes_4_7_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_5_6), //i
    .io_resetPartialC        (io_resetPartialC_5_6       ), //i
    .io_outputA              (pes_5_6_io_outputA[7:0]    ), //o
    .io_outputB              (pes_5_6_io_outputB[7:0]    ), //o
    .io_outputC              (pes_5_6_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_5_7 (
    .io_inputA               (pes_5_6_io_outputA[7:0]    ), //i
    .io_inputB               (pes_4_7_io_outputB[7:0]    ), //i
    .io_inputC               (pes_4_8_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_5_7), //i
    .io_resetPartialC        (io_resetPartialC_5_7       ), //i
    .io_outputA              (pes_5_7_io_outputA[7:0]    ), //o
    .io_outputB              (pes_5_7_io_outputB[7:0]    ), //o
    .io_outputC              (pes_5_7_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_5_8 (
    .io_inputA               (pes_5_7_io_outputA[7:0]    ), //i
    .io_inputB               (pes_4_8_io_outputB[7:0]    ), //i
    .io_inputC               (pes_4_9_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_5_8), //i
    .io_resetPartialC        (io_resetPartialC_5_8       ), //i
    .io_outputA              (pes_5_8_io_outputA[7:0]    ), //o
    .io_outputB              (pes_5_8_io_outputB[7:0]    ), //o
    .io_outputC              (pes_5_8_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_5_9 (
    .io_inputA               (pes_5_8_io_outputA[7:0]    ), //i
    .io_inputB               (pes_4_9_io_outputB[7:0]    ), //i
    .io_inputC               (pes_4_10_io_outputC[25:0]  ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_5_9), //i
    .io_resetPartialC        (io_resetPartialC_5_9       ), //i
    .io_outputA              (pes_5_9_io_outputA[7:0]    ), //o
    .io_outputB              (pes_5_9_io_outputB[7:0]    ), //o
    .io_outputC              (pes_5_9_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_5_10 (
    .io_inputA               (pes_5_9_io_outputA[7:0]     ), //i
    .io_inputB               (pes_4_10_io_outputB[7:0]    ), //i
    .io_inputC               (pes_4_11_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_5_10), //i
    .io_resetPartialC        (io_resetPartialC_5_10       ), //i
    .io_outputA              (pes_5_10_io_outputA[7:0]    ), //o
    .io_outputB              (pes_5_10_io_outputB[7:0]    ), //o
    .io_outputC              (pes_5_10_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_5_11 (
    .io_inputA               (pes_5_10_io_outputA[7:0]    ), //i
    .io_inputB               (pes_4_11_io_outputB[7:0]    ), //i
    .io_inputC               (pes_4_12_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_5_11), //i
    .io_resetPartialC        (io_resetPartialC_5_11       ), //i
    .io_outputA              (pes_5_11_io_outputA[7:0]    ), //o
    .io_outputB              (pes_5_11_io_outputB[7:0]    ), //o
    .io_outputC              (pes_5_11_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_5_12 (
    .io_inputA               (pes_5_11_io_outputA[7:0]    ), //i
    .io_inputB               (pes_4_12_io_outputB[7:0]    ), //i
    .io_inputC               (pes_4_13_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_5_12), //i
    .io_resetPartialC        (io_resetPartialC_5_12       ), //i
    .io_outputA              (pes_5_12_io_outputA[7:0]    ), //o
    .io_outputB              (pes_5_12_io_outputB[7:0]    ), //o
    .io_outputC              (pes_5_12_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_5_13 (
    .io_inputA               (pes_5_12_io_outputA[7:0]    ), //i
    .io_inputB               (pes_4_13_io_outputB[7:0]    ), //i
    .io_inputC               (pes_4_14_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_5_13), //i
    .io_resetPartialC        (io_resetPartialC_5_13       ), //i
    .io_outputA              (pes_5_13_io_outputA[7:0]    ), //o
    .io_outputB              (pes_5_13_io_outputB[7:0]    ), //o
    .io_outputC              (pes_5_13_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_5_14 (
    .io_inputA               (pes_5_13_io_outputA[7:0]    ), //i
    .io_inputB               (pes_4_14_io_outputB[7:0]    ), //i
    .io_inputC               (pes_4_15_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_5_14), //i
    .io_resetPartialC        (io_resetPartialC_5_14       ), //i
    .io_outputA              (pes_5_14_io_outputA[7:0]    ), //o
    .io_outputB              (pes_5_14_io_outputB[7:0]    ), //o
    .io_outputC              (pes_5_14_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_15 pes_5_15 (
    .io_inputA               (pes_5_14_io_outputA[7:0]    ), //i
    .io_inputB               (pes_4_15_io_outputB[7:0]    ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_5_15), //i
    .io_resetPartialC        (io_resetPartialC_5_15       ), //i
    .io_outputB              (pes_5_15_io_outputB[7:0]    ), //o
    .io_outputC              (pes_5_15_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_6_0 (
    .io_inputA               (skewBuffer_io_output_6[7:0]), //i
    .io_inputB               (pes_5_0_io_outputB[7:0]    ), //i
    .io_inputC               (pes_5_1_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_6_0), //i
    .io_resetPartialC        (io_resetPartialC_6_0       ), //i
    .io_outputA              (pes_6_0_io_outputA[7:0]    ), //o
    .io_outputB              (pes_6_0_io_outputB[7:0]    ), //o
    .io_outputC              (pes_6_0_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_6_1 (
    .io_inputA               (pes_6_0_io_outputA[7:0]    ), //i
    .io_inputB               (pes_5_1_io_outputB[7:0]    ), //i
    .io_inputC               (pes_5_2_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_6_1), //i
    .io_resetPartialC        (io_resetPartialC_6_1       ), //i
    .io_outputA              (pes_6_1_io_outputA[7:0]    ), //o
    .io_outputB              (pes_6_1_io_outputB[7:0]    ), //o
    .io_outputC              (pes_6_1_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_6_2 (
    .io_inputA               (pes_6_1_io_outputA[7:0]    ), //i
    .io_inputB               (pes_5_2_io_outputB[7:0]    ), //i
    .io_inputC               (pes_5_3_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_6_2), //i
    .io_resetPartialC        (io_resetPartialC_6_2       ), //i
    .io_outputA              (pes_6_2_io_outputA[7:0]    ), //o
    .io_outputB              (pes_6_2_io_outputB[7:0]    ), //o
    .io_outputC              (pes_6_2_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_6_3 (
    .io_inputA               (pes_6_2_io_outputA[7:0]    ), //i
    .io_inputB               (pes_5_3_io_outputB[7:0]    ), //i
    .io_inputC               (pes_5_4_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_6_3), //i
    .io_resetPartialC        (io_resetPartialC_6_3       ), //i
    .io_outputA              (pes_6_3_io_outputA[7:0]    ), //o
    .io_outputB              (pes_6_3_io_outputB[7:0]    ), //o
    .io_outputC              (pes_6_3_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_6_4 (
    .io_inputA               (pes_6_3_io_outputA[7:0]    ), //i
    .io_inputB               (pes_5_4_io_outputB[7:0]    ), //i
    .io_inputC               (pes_5_5_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_6_4), //i
    .io_resetPartialC        (io_resetPartialC_6_4       ), //i
    .io_outputA              (pes_6_4_io_outputA[7:0]    ), //o
    .io_outputB              (pes_6_4_io_outputB[7:0]    ), //o
    .io_outputC              (pes_6_4_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_6_5 (
    .io_inputA               (pes_6_4_io_outputA[7:0]    ), //i
    .io_inputB               (pes_5_5_io_outputB[7:0]    ), //i
    .io_inputC               (pes_5_6_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_6_5), //i
    .io_resetPartialC        (io_resetPartialC_6_5       ), //i
    .io_outputA              (pes_6_5_io_outputA[7:0]    ), //o
    .io_outputB              (pes_6_5_io_outputB[7:0]    ), //o
    .io_outputC              (pes_6_5_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_6_6 (
    .io_inputA               (pes_6_5_io_outputA[7:0]    ), //i
    .io_inputB               (pes_5_6_io_outputB[7:0]    ), //i
    .io_inputC               (pes_5_7_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_6_6), //i
    .io_resetPartialC        (io_resetPartialC_6_6       ), //i
    .io_outputA              (pes_6_6_io_outputA[7:0]    ), //o
    .io_outputB              (pes_6_6_io_outputB[7:0]    ), //o
    .io_outputC              (pes_6_6_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_6_7 (
    .io_inputA               (pes_6_6_io_outputA[7:0]    ), //i
    .io_inputB               (pes_5_7_io_outputB[7:0]    ), //i
    .io_inputC               (pes_5_8_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_6_7), //i
    .io_resetPartialC        (io_resetPartialC_6_7       ), //i
    .io_outputA              (pes_6_7_io_outputA[7:0]    ), //o
    .io_outputB              (pes_6_7_io_outputB[7:0]    ), //o
    .io_outputC              (pes_6_7_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_6_8 (
    .io_inputA               (pes_6_7_io_outputA[7:0]    ), //i
    .io_inputB               (pes_5_8_io_outputB[7:0]    ), //i
    .io_inputC               (pes_5_9_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_6_8), //i
    .io_resetPartialC        (io_resetPartialC_6_8       ), //i
    .io_outputA              (pes_6_8_io_outputA[7:0]    ), //o
    .io_outputB              (pes_6_8_io_outputB[7:0]    ), //o
    .io_outputC              (pes_6_8_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_6_9 (
    .io_inputA               (pes_6_8_io_outputA[7:0]    ), //i
    .io_inputB               (pes_5_9_io_outputB[7:0]    ), //i
    .io_inputC               (pes_5_10_io_outputC[25:0]  ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_6_9), //i
    .io_resetPartialC        (io_resetPartialC_6_9       ), //i
    .io_outputA              (pes_6_9_io_outputA[7:0]    ), //o
    .io_outputB              (pes_6_9_io_outputB[7:0]    ), //o
    .io_outputC              (pes_6_9_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_6_10 (
    .io_inputA               (pes_6_9_io_outputA[7:0]     ), //i
    .io_inputB               (pes_5_10_io_outputB[7:0]    ), //i
    .io_inputC               (pes_5_11_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_6_10), //i
    .io_resetPartialC        (io_resetPartialC_6_10       ), //i
    .io_outputA              (pes_6_10_io_outputA[7:0]    ), //o
    .io_outputB              (pes_6_10_io_outputB[7:0]    ), //o
    .io_outputC              (pes_6_10_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_6_11 (
    .io_inputA               (pes_6_10_io_outputA[7:0]    ), //i
    .io_inputB               (pes_5_11_io_outputB[7:0]    ), //i
    .io_inputC               (pes_5_12_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_6_11), //i
    .io_resetPartialC        (io_resetPartialC_6_11       ), //i
    .io_outputA              (pes_6_11_io_outputA[7:0]    ), //o
    .io_outputB              (pes_6_11_io_outputB[7:0]    ), //o
    .io_outputC              (pes_6_11_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_6_12 (
    .io_inputA               (pes_6_11_io_outputA[7:0]    ), //i
    .io_inputB               (pes_5_12_io_outputB[7:0]    ), //i
    .io_inputC               (pes_5_13_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_6_12), //i
    .io_resetPartialC        (io_resetPartialC_6_12       ), //i
    .io_outputA              (pes_6_12_io_outputA[7:0]    ), //o
    .io_outputB              (pes_6_12_io_outputB[7:0]    ), //o
    .io_outputC              (pes_6_12_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_6_13 (
    .io_inputA               (pes_6_12_io_outputA[7:0]    ), //i
    .io_inputB               (pes_5_13_io_outputB[7:0]    ), //i
    .io_inputC               (pes_5_14_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_6_13), //i
    .io_resetPartialC        (io_resetPartialC_6_13       ), //i
    .io_outputA              (pes_6_13_io_outputA[7:0]    ), //o
    .io_outputB              (pes_6_13_io_outputB[7:0]    ), //o
    .io_outputC              (pes_6_13_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_6_14 (
    .io_inputA               (pes_6_13_io_outputA[7:0]    ), //i
    .io_inputB               (pes_5_14_io_outputB[7:0]    ), //i
    .io_inputC               (pes_5_15_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_6_14), //i
    .io_resetPartialC        (io_resetPartialC_6_14       ), //i
    .io_outputA              (pes_6_14_io_outputA[7:0]    ), //o
    .io_outputB              (pes_6_14_io_outputB[7:0]    ), //o
    .io_outputC              (pes_6_14_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_15 pes_6_15 (
    .io_inputA               (pes_6_14_io_outputA[7:0]    ), //i
    .io_inputB               (pes_5_15_io_outputB[7:0]    ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_6_15), //i
    .io_resetPartialC        (io_resetPartialC_6_15       ), //i
    .io_outputB              (pes_6_15_io_outputB[7:0]    ), //o
    .io_outputC              (pes_6_15_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_7_0 (
    .io_inputA               (skewBuffer_io_output_7[7:0]), //i
    .io_inputB               (pes_6_0_io_outputB[7:0]    ), //i
    .io_inputC               (pes_6_1_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_7_0), //i
    .io_resetPartialC        (io_resetPartialC_7_0       ), //i
    .io_outputA              (pes_7_0_io_outputA[7:0]    ), //o
    .io_outputB              (pes_7_0_io_outputB[7:0]    ), //o
    .io_outputC              (pes_7_0_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_7_1 (
    .io_inputA               (pes_7_0_io_outputA[7:0]    ), //i
    .io_inputB               (pes_6_1_io_outputB[7:0]    ), //i
    .io_inputC               (pes_6_2_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_7_1), //i
    .io_resetPartialC        (io_resetPartialC_7_1       ), //i
    .io_outputA              (pes_7_1_io_outputA[7:0]    ), //o
    .io_outputB              (pes_7_1_io_outputB[7:0]    ), //o
    .io_outputC              (pes_7_1_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_7_2 (
    .io_inputA               (pes_7_1_io_outputA[7:0]    ), //i
    .io_inputB               (pes_6_2_io_outputB[7:0]    ), //i
    .io_inputC               (pes_6_3_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_7_2), //i
    .io_resetPartialC        (io_resetPartialC_7_2       ), //i
    .io_outputA              (pes_7_2_io_outputA[7:0]    ), //o
    .io_outputB              (pes_7_2_io_outputB[7:0]    ), //o
    .io_outputC              (pes_7_2_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_7_3 (
    .io_inputA               (pes_7_2_io_outputA[7:0]    ), //i
    .io_inputB               (pes_6_3_io_outputB[7:0]    ), //i
    .io_inputC               (pes_6_4_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_7_3), //i
    .io_resetPartialC        (io_resetPartialC_7_3       ), //i
    .io_outputA              (pes_7_3_io_outputA[7:0]    ), //o
    .io_outputB              (pes_7_3_io_outputB[7:0]    ), //o
    .io_outputC              (pes_7_3_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_7_4 (
    .io_inputA               (pes_7_3_io_outputA[7:0]    ), //i
    .io_inputB               (pes_6_4_io_outputB[7:0]    ), //i
    .io_inputC               (pes_6_5_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_7_4), //i
    .io_resetPartialC        (io_resetPartialC_7_4       ), //i
    .io_outputA              (pes_7_4_io_outputA[7:0]    ), //o
    .io_outputB              (pes_7_4_io_outputB[7:0]    ), //o
    .io_outputC              (pes_7_4_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_7_5 (
    .io_inputA               (pes_7_4_io_outputA[7:0]    ), //i
    .io_inputB               (pes_6_5_io_outputB[7:0]    ), //i
    .io_inputC               (pes_6_6_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_7_5), //i
    .io_resetPartialC        (io_resetPartialC_7_5       ), //i
    .io_outputA              (pes_7_5_io_outputA[7:0]    ), //o
    .io_outputB              (pes_7_5_io_outputB[7:0]    ), //o
    .io_outputC              (pes_7_5_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_7_6 (
    .io_inputA               (pes_7_5_io_outputA[7:0]    ), //i
    .io_inputB               (pes_6_6_io_outputB[7:0]    ), //i
    .io_inputC               (pes_6_7_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_7_6), //i
    .io_resetPartialC        (io_resetPartialC_7_6       ), //i
    .io_outputA              (pes_7_6_io_outputA[7:0]    ), //o
    .io_outputB              (pes_7_6_io_outputB[7:0]    ), //o
    .io_outputC              (pes_7_6_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_7_7 (
    .io_inputA               (pes_7_6_io_outputA[7:0]    ), //i
    .io_inputB               (pes_6_7_io_outputB[7:0]    ), //i
    .io_inputC               (pes_6_8_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_7_7), //i
    .io_resetPartialC        (io_resetPartialC_7_7       ), //i
    .io_outputA              (pes_7_7_io_outputA[7:0]    ), //o
    .io_outputB              (pes_7_7_io_outputB[7:0]    ), //o
    .io_outputC              (pes_7_7_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_7_8 (
    .io_inputA               (pes_7_7_io_outputA[7:0]    ), //i
    .io_inputB               (pes_6_8_io_outputB[7:0]    ), //i
    .io_inputC               (pes_6_9_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_7_8), //i
    .io_resetPartialC        (io_resetPartialC_7_8       ), //i
    .io_outputA              (pes_7_8_io_outputA[7:0]    ), //o
    .io_outputB              (pes_7_8_io_outputB[7:0]    ), //o
    .io_outputC              (pes_7_8_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_7_9 (
    .io_inputA               (pes_7_8_io_outputA[7:0]    ), //i
    .io_inputB               (pes_6_9_io_outputB[7:0]    ), //i
    .io_inputC               (pes_6_10_io_outputC[25:0]  ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_7_9), //i
    .io_resetPartialC        (io_resetPartialC_7_9       ), //i
    .io_outputA              (pes_7_9_io_outputA[7:0]    ), //o
    .io_outputB              (pes_7_9_io_outputB[7:0]    ), //o
    .io_outputC              (pes_7_9_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_7_10 (
    .io_inputA               (pes_7_9_io_outputA[7:0]     ), //i
    .io_inputB               (pes_6_10_io_outputB[7:0]    ), //i
    .io_inputC               (pes_6_11_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_7_10), //i
    .io_resetPartialC        (io_resetPartialC_7_10       ), //i
    .io_outputA              (pes_7_10_io_outputA[7:0]    ), //o
    .io_outputB              (pes_7_10_io_outputB[7:0]    ), //o
    .io_outputC              (pes_7_10_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_7_11 (
    .io_inputA               (pes_7_10_io_outputA[7:0]    ), //i
    .io_inputB               (pes_6_11_io_outputB[7:0]    ), //i
    .io_inputC               (pes_6_12_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_7_11), //i
    .io_resetPartialC        (io_resetPartialC_7_11       ), //i
    .io_outputA              (pes_7_11_io_outputA[7:0]    ), //o
    .io_outputB              (pes_7_11_io_outputB[7:0]    ), //o
    .io_outputC              (pes_7_11_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_7_12 (
    .io_inputA               (pes_7_11_io_outputA[7:0]    ), //i
    .io_inputB               (pes_6_12_io_outputB[7:0]    ), //i
    .io_inputC               (pes_6_13_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_7_12), //i
    .io_resetPartialC        (io_resetPartialC_7_12       ), //i
    .io_outputA              (pes_7_12_io_outputA[7:0]    ), //o
    .io_outputB              (pes_7_12_io_outputB[7:0]    ), //o
    .io_outputC              (pes_7_12_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_7_13 (
    .io_inputA               (pes_7_12_io_outputA[7:0]    ), //i
    .io_inputB               (pes_6_13_io_outputB[7:0]    ), //i
    .io_inputC               (pes_6_14_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_7_13), //i
    .io_resetPartialC        (io_resetPartialC_7_13       ), //i
    .io_outputA              (pes_7_13_io_outputA[7:0]    ), //o
    .io_outputB              (pes_7_13_io_outputB[7:0]    ), //o
    .io_outputC              (pes_7_13_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_7_14 (
    .io_inputA               (pes_7_13_io_outputA[7:0]    ), //i
    .io_inputB               (pes_6_14_io_outputB[7:0]    ), //i
    .io_inputC               (pes_6_15_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_7_14), //i
    .io_resetPartialC        (io_resetPartialC_7_14       ), //i
    .io_outputA              (pes_7_14_io_outputA[7:0]    ), //o
    .io_outputB              (pes_7_14_io_outputB[7:0]    ), //o
    .io_outputC              (pes_7_14_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_15 pes_7_15 (
    .io_inputA               (pes_7_14_io_outputA[7:0]    ), //i
    .io_inputB               (pes_6_15_io_outputB[7:0]    ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_7_15), //i
    .io_resetPartialC        (io_resetPartialC_7_15       ), //i
    .io_outputB              (pes_7_15_io_outputB[7:0]    ), //o
    .io_outputC              (pes_7_15_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_8_0 (
    .io_inputA               (skewBuffer_io_output_8[7:0]), //i
    .io_inputB               (pes_7_0_io_outputB[7:0]    ), //i
    .io_inputC               (pes_7_1_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_8_0), //i
    .io_resetPartialC        (io_resetPartialC_8_0       ), //i
    .io_outputA              (pes_8_0_io_outputA[7:0]    ), //o
    .io_outputB              (pes_8_0_io_outputB[7:0]    ), //o
    .io_outputC              (pes_8_0_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_8_1 (
    .io_inputA               (pes_8_0_io_outputA[7:0]    ), //i
    .io_inputB               (pes_7_1_io_outputB[7:0]    ), //i
    .io_inputC               (pes_7_2_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_8_1), //i
    .io_resetPartialC        (io_resetPartialC_8_1       ), //i
    .io_outputA              (pes_8_1_io_outputA[7:0]    ), //o
    .io_outputB              (pes_8_1_io_outputB[7:0]    ), //o
    .io_outputC              (pes_8_1_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_8_2 (
    .io_inputA               (pes_8_1_io_outputA[7:0]    ), //i
    .io_inputB               (pes_7_2_io_outputB[7:0]    ), //i
    .io_inputC               (pes_7_3_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_8_2), //i
    .io_resetPartialC        (io_resetPartialC_8_2       ), //i
    .io_outputA              (pes_8_2_io_outputA[7:0]    ), //o
    .io_outputB              (pes_8_2_io_outputB[7:0]    ), //o
    .io_outputC              (pes_8_2_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_8_3 (
    .io_inputA               (pes_8_2_io_outputA[7:0]    ), //i
    .io_inputB               (pes_7_3_io_outputB[7:0]    ), //i
    .io_inputC               (pes_7_4_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_8_3), //i
    .io_resetPartialC        (io_resetPartialC_8_3       ), //i
    .io_outputA              (pes_8_3_io_outputA[7:0]    ), //o
    .io_outputB              (pes_8_3_io_outputB[7:0]    ), //o
    .io_outputC              (pes_8_3_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_8_4 (
    .io_inputA               (pes_8_3_io_outputA[7:0]    ), //i
    .io_inputB               (pes_7_4_io_outputB[7:0]    ), //i
    .io_inputC               (pes_7_5_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_8_4), //i
    .io_resetPartialC        (io_resetPartialC_8_4       ), //i
    .io_outputA              (pes_8_4_io_outputA[7:0]    ), //o
    .io_outputB              (pes_8_4_io_outputB[7:0]    ), //o
    .io_outputC              (pes_8_4_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_8_5 (
    .io_inputA               (pes_8_4_io_outputA[7:0]    ), //i
    .io_inputB               (pes_7_5_io_outputB[7:0]    ), //i
    .io_inputC               (pes_7_6_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_8_5), //i
    .io_resetPartialC        (io_resetPartialC_8_5       ), //i
    .io_outputA              (pes_8_5_io_outputA[7:0]    ), //o
    .io_outputB              (pes_8_5_io_outputB[7:0]    ), //o
    .io_outputC              (pes_8_5_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_8_6 (
    .io_inputA               (pes_8_5_io_outputA[7:0]    ), //i
    .io_inputB               (pes_7_6_io_outputB[7:0]    ), //i
    .io_inputC               (pes_7_7_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_8_6), //i
    .io_resetPartialC        (io_resetPartialC_8_6       ), //i
    .io_outputA              (pes_8_6_io_outputA[7:0]    ), //o
    .io_outputB              (pes_8_6_io_outputB[7:0]    ), //o
    .io_outputC              (pes_8_6_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_8_7 (
    .io_inputA               (pes_8_6_io_outputA[7:0]    ), //i
    .io_inputB               (pes_7_7_io_outputB[7:0]    ), //i
    .io_inputC               (pes_7_8_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_8_7), //i
    .io_resetPartialC        (io_resetPartialC_8_7       ), //i
    .io_outputA              (pes_8_7_io_outputA[7:0]    ), //o
    .io_outputB              (pes_8_7_io_outputB[7:0]    ), //o
    .io_outputC              (pes_8_7_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_8_8 (
    .io_inputA               (pes_8_7_io_outputA[7:0]    ), //i
    .io_inputB               (pes_7_8_io_outputB[7:0]    ), //i
    .io_inputC               (pes_7_9_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_8_8), //i
    .io_resetPartialC        (io_resetPartialC_8_8       ), //i
    .io_outputA              (pes_8_8_io_outputA[7:0]    ), //o
    .io_outputB              (pes_8_8_io_outputB[7:0]    ), //o
    .io_outputC              (pes_8_8_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_8_9 (
    .io_inputA               (pes_8_8_io_outputA[7:0]    ), //i
    .io_inputB               (pes_7_9_io_outputB[7:0]    ), //i
    .io_inputC               (pes_7_10_io_outputC[25:0]  ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_8_9), //i
    .io_resetPartialC        (io_resetPartialC_8_9       ), //i
    .io_outputA              (pes_8_9_io_outputA[7:0]    ), //o
    .io_outputB              (pes_8_9_io_outputB[7:0]    ), //o
    .io_outputC              (pes_8_9_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_8_10 (
    .io_inputA               (pes_8_9_io_outputA[7:0]     ), //i
    .io_inputB               (pes_7_10_io_outputB[7:0]    ), //i
    .io_inputC               (pes_7_11_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_8_10), //i
    .io_resetPartialC        (io_resetPartialC_8_10       ), //i
    .io_outputA              (pes_8_10_io_outputA[7:0]    ), //o
    .io_outputB              (pes_8_10_io_outputB[7:0]    ), //o
    .io_outputC              (pes_8_10_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_8_11 (
    .io_inputA               (pes_8_10_io_outputA[7:0]    ), //i
    .io_inputB               (pes_7_11_io_outputB[7:0]    ), //i
    .io_inputC               (pes_7_12_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_8_11), //i
    .io_resetPartialC        (io_resetPartialC_8_11       ), //i
    .io_outputA              (pes_8_11_io_outputA[7:0]    ), //o
    .io_outputB              (pes_8_11_io_outputB[7:0]    ), //o
    .io_outputC              (pes_8_11_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_8_12 (
    .io_inputA               (pes_8_11_io_outputA[7:0]    ), //i
    .io_inputB               (pes_7_12_io_outputB[7:0]    ), //i
    .io_inputC               (pes_7_13_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_8_12), //i
    .io_resetPartialC        (io_resetPartialC_8_12       ), //i
    .io_outputA              (pes_8_12_io_outputA[7:0]    ), //o
    .io_outputB              (pes_8_12_io_outputB[7:0]    ), //o
    .io_outputC              (pes_8_12_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_8_13 (
    .io_inputA               (pes_8_12_io_outputA[7:0]    ), //i
    .io_inputB               (pes_7_13_io_outputB[7:0]    ), //i
    .io_inputC               (pes_7_14_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_8_13), //i
    .io_resetPartialC        (io_resetPartialC_8_13       ), //i
    .io_outputA              (pes_8_13_io_outputA[7:0]    ), //o
    .io_outputB              (pes_8_13_io_outputB[7:0]    ), //o
    .io_outputC              (pes_8_13_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_8_14 (
    .io_inputA               (pes_8_13_io_outputA[7:0]    ), //i
    .io_inputB               (pes_7_14_io_outputB[7:0]    ), //i
    .io_inputC               (pes_7_15_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_8_14), //i
    .io_resetPartialC        (io_resetPartialC_8_14       ), //i
    .io_outputA              (pes_8_14_io_outputA[7:0]    ), //o
    .io_outputB              (pes_8_14_io_outputB[7:0]    ), //o
    .io_outputC              (pes_8_14_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_15 pes_8_15 (
    .io_inputA               (pes_8_14_io_outputA[7:0]    ), //i
    .io_inputB               (pes_7_15_io_outputB[7:0]    ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_8_15), //i
    .io_resetPartialC        (io_resetPartialC_8_15       ), //i
    .io_outputB              (pes_8_15_io_outputB[7:0]    ), //o
    .io_outputC              (pes_8_15_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_9_0 (
    .io_inputA               (skewBuffer_io_output_9[7:0]), //i
    .io_inputB               (pes_8_0_io_outputB[7:0]    ), //i
    .io_inputC               (pes_8_1_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_9_0), //i
    .io_resetPartialC        (io_resetPartialC_9_0       ), //i
    .io_outputA              (pes_9_0_io_outputA[7:0]    ), //o
    .io_outputB              (pes_9_0_io_outputB[7:0]    ), //o
    .io_outputC              (pes_9_0_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_9_1 (
    .io_inputA               (pes_9_0_io_outputA[7:0]    ), //i
    .io_inputB               (pes_8_1_io_outputB[7:0]    ), //i
    .io_inputC               (pes_8_2_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_9_1), //i
    .io_resetPartialC        (io_resetPartialC_9_1       ), //i
    .io_outputA              (pes_9_1_io_outputA[7:0]    ), //o
    .io_outputB              (pes_9_1_io_outputB[7:0]    ), //o
    .io_outputC              (pes_9_1_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_9_2 (
    .io_inputA               (pes_9_1_io_outputA[7:0]    ), //i
    .io_inputB               (pes_8_2_io_outputB[7:0]    ), //i
    .io_inputC               (pes_8_3_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_9_2), //i
    .io_resetPartialC        (io_resetPartialC_9_2       ), //i
    .io_outputA              (pes_9_2_io_outputA[7:0]    ), //o
    .io_outputB              (pes_9_2_io_outputB[7:0]    ), //o
    .io_outputC              (pes_9_2_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_9_3 (
    .io_inputA               (pes_9_2_io_outputA[7:0]    ), //i
    .io_inputB               (pes_8_3_io_outputB[7:0]    ), //i
    .io_inputC               (pes_8_4_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_9_3), //i
    .io_resetPartialC        (io_resetPartialC_9_3       ), //i
    .io_outputA              (pes_9_3_io_outputA[7:0]    ), //o
    .io_outputB              (pes_9_3_io_outputB[7:0]    ), //o
    .io_outputC              (pes_9_3_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_9_4 (
    .io_inputA               (pes_9_3_io_outputA[7:0]    ), //i
    .io_inputB               (pes_8_4_io_outputB[7:0]    ), //i
    .io_inputC               (pes_8_5_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_9_4), //i
    .io_resetPartialC        (io_resetPartialC_9_4       ), //i
    .io_outputA              (pes_9_4_io_outputA[7:0]    ), //o
    .io_outputB              (pes_9_4_io_outputB[7:0]    ), //o
    .io_outputC              (pes_9_4_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_9_5 (
    .io_inputA               (pes_9_4_io_outputA[7:0]    ), //i
    .io_inputB               (pes_8_5_io_outputB[7:0]    ), //i
    .io_inputC               (pes_8_6_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_9_5), //i
    .io_resetPartialC        (io_resetPartialC_9_5       ), //i
    .io_outputA              (pes_9_5_io_outputA[7:0]    ), //o
    .io_outputB              (pes_9_5_io_outputB[7:0]    ), //o
    .io_outputC              (pes_9_5_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_9_6 (
    .io_inputA               (pes_9_5_io_outputA[7:0]    ), //i
    .io_inputB               (pes_8_6_io_outputB[7:0]    ), //i
    .io_inputC               (pes_8_7_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_9_6), //i
    .io_resetPartialC        (io_resetPartialC_9_6       ), //i
    .io_outputA              (pes_9_6_io_outputA[7:0]    ), //o
    .io_outputB              (pes_9_6_io_outputB[7:0]    ), //o
    .io_outputC              (pes_9_6_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_9_7 (
    .io_inputA               (pes_9_6_io_outputA[7:0]    ), //i
    .io_inputB               (pes_8_7_io_outputB[7:0]    ), //i
    .io_inputC               (pes_8_8_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_9_7), //i
    .io_resetPartialC        (io_resetPartialC_9_7       ), //i
    .io_outputA              (pes_9_7_io_outputA[7:0]    ), //o
    .io_outputB              (pes_9_7_io_outputB[7:0]    ), //o
    .io_outputC              (pes_9_7_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_9_8 (
    .io_inputA               (pes_9_7_io_outputA[7:0]    ), //i
    .io_inputB               (pes_8_8_io_outputB[7:0]    ), //i
    .io_inputC               (pes_8_9_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_9_8), //i
    .io_resetPartialC        (io_resetPartialC_9_8       ), //i
    .io_outputA              (pes_9_8_io_outputA[7:0]    ), //o
    .io_outputB              (pes_9_8_io_outputB[7:0]    ), //o
    .io_outputC              (pes_9_8_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_9_9 (
    .io_inputA               (pes_9_8_io_outputA[7:0]    ), //i
    .io_inputB               (pes_8_9_io_outputB[7:0]    ), //i
    .io_inputC               (pes_8_10_io_outputC[25:0]  ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_9_9), //i
    .io_resetPartialC        (io_resetPartialC_9_9       ), //i
    .io_outputA              (pes_9_9_io_outputA[7:0]    ), //o
    .io_outputB              (pes_9_9_io_outputB[7:0]    ), //o
    .io_outputC              (pes_9_9_io_outputC[25:0]   ), //o
    .clk                     (clk                        ), //i
    .reset                   (reset                      )  //i
  );
  ProcessingElement_16 pes_9_10 (
    .io_inputA               (pes_9_9_io_outputA[7:0]     ), //i
    .io_inputB               (pes_8_10_io_outputB[7:0]    ), //i
    .io_inputC               (pes_8_11_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_9_10), //i
    .io_resetPartialC        (io_resetPartialC_9_10       ), //i
    .io_outputA              (pes_9_10_io_outputA[7:0]    ), //o
    .io_outputB              (pes_9_10_io_outputB[7:0]    ), //o
    .io_outputC              (pes_9_10_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_9_11 (
    .io_inputA               (pes_9_10_io_outputA[7:0]    ), //i
    .io_inputB               (pes_8_11_io_outputB[7:0]    ), //i
    .io_inputC               (pes_8_12_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_9_11), //i
    .io_resetPartialC        (io_resetPartialC_9_11       ), //i
    .io_outputA              (pes_9_11_io_outputA[7:0]    ), //o
    .io_outputB              (pes_9_11_io_outputB[7:0]    ), //o
    .io_outputC              (pes_9_11_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_9_12 (
    .io_inputA               (pes_9_11_io_outputA[7:0]    ), //i
    .io_inputB               (pes_8_12_io_outputB[7:0]    ), //i
    .io_inputC               (pes_8_13_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_9_12), //i
    .io_resetPartialC        (io_resetPartialC_9_12       ), //i
    .io_outputA              (pes_9_12_io_outputA[7:0]    ), //o
    .io_outputB              (pes_9_12_io_outputB[7:0]    ), //o
    .io_outputC              (pes_9_12_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_9_13 (
    .io_inputA               (pes_9_12_io_outputA[7:0]    ), //i
    .io_inputB               (pes_8_13_io_outputB[7:0]    ), //i
    .io_inputC               (pes_8_14_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_9_13), //i
    .io_resetPartialC        (io_resetPartialC_9_13       ), //i
    .io_outputA              (pes_9_13_io_outputA[7:0]    ), //o
    .io_outputB              (pes_9_13_io_outputB[7:0]    ), //o
    .io_outputC              (pes_9_13_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_9_14 (
    .io_inputA               (pes_9_13_io_outputA[7:0]    ), //i
    .io_inputB               (pes_8_14_io_outputB[7:0]    ), //i
    .io_inputC               (pes_8_15_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_9_14), //i
    .io_resetPartialC        (io_resetPartialC_9_14       ), //i
    .io_outputA              (pes_9_14_io_outputA[7:0]    ), //o
    .io_outputB              (pes_9_14_io_outputB[7:0]    ), //o
    .io_outputC              (pes_9_14_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_15 pes_9_15 (
    .io_inputA               (pes_9_14_io_outputA[7:0]    ), //i
    .io_inputB               (pes_8_15_io_outputB[7:0]    ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_9_15), //i
    .io_resetPartialC        (io_resetPartialC_9_15       ), //i
    .io_outputB              (pes_9_15_io_outputB[7:0]    ), //o
    .io_outputC              (pes_9_15_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_10_0 (
    .io_inputA               (skewBuffer_io_output_10[7:0]), //i
    .io_inputB               (pes_9_0_io_outputB[7:0]     ), //i
    .io_inputC               (pes_9_1_io_outputC[25:0]    ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_10_0), //i
    .io_resetPartialC        (io_resetPartialC_10_0       ), //i
    .io_outputA              (pes_10_0_io_outputA[7:0]    ), //o
    .io_outputB              (pes_10_0_io_outputB[7:0]    ), //o
    .io_outputC              (pes_10_0_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_10_1 (
    .io_inputA               (pes_10_0_io_outputA[7:0]    ), //i
    .io_inputB               (pes_9_1_io_outputB[7:0]     ), //i
    .io_inputC               (pes_9_2_io_outputC[25:0]    ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_10_1), //i
    .io_resetPartialC        (io_resetPartialC_10_1       ), //i
    .io_outputA              (pes_10_1_io_outputA[7:0]    ), //o
    .io_outputB              (pes_10_1_io_outputB[7:0]    ), //o
    .io_outputC              (pes_10_1_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_10_2 (
    .io_inputA               (pes_10_1_io_outputA[7:0]    ), //i
    .io_inputB               (pes_9_2_io_outputB[7:0]     ), //i
    .io_inputC               (pes_9_3_io_outputC[25:0]    ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_10_2), //i
    .io_resetPartialC        (io_resetPartialC_10_2       ), //i
    .io_outputA              (pes_10_2_io_outputA[7:0]    ), //o
    .io_outputB              (pes_10_2_io_outputB[7:0]    ), //o
    .io_outputC              (pes_10_2_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_10_3 (
    .io_inputA               (pes_10_2_io_outputA[7:0]    ), //i
    .io_inputB               (pes_9_3_io_outputB[7:0]     ), //i
    .io_inputC               (pes_9_4_io_outputC[25:0]    ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_10_3), //i
    .io_resetPartialC        (io_resetPartialC_10_3       ), //i
    .io_outputA              (pes_10_3_io_outputA[7:0]    ), //o
    .io_outputB              (pes_10_3_io_outputB[7:0]    ), //o
    .io_outputC              (pes_10_3_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_10_4 (
    .io_inputA               (pes_10_3_io_outputA[7:0]    ), //i
    .io_inputB               (pes_9_4_io_outputB[7:0]     ), //i
    .io_inputC               (pes_9_5_io_outputC[25:0]    ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_10_4), //i
    .io_resetPartialC        (io_resetPartialC_10_4       ), //i
    .io_outputA              (pes_10_4_io_outputA[7:0]    ), //o
    .io_outputB              (pes_10_4_io_outputB[7:0]    ), //o
    .io_outputC              (pes_10_4_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_10_5 (
    .io_inputA               (pes_10_4_io_outputA[7:0]    ), //i
    .io_inputB               (pes_9_5_io_outputB[7:0]     ), //i
    .io_inputC               (pes_9_6_io_outputC[25:0]    ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_10_5), //i
    .io_resetPartialC        (io_resetPartialC_10_5       ), //i
    .io_outputA              (pes_10_5_io_outputA[7:0]    ), //o
    .io_outputB              (pes_10_5_io_outputB[7:0]    ), //o
    .io_outputC              (pes_10_5_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_10_6 (
    .io_inputA               (pes_10_5_io_outputA[7:0]    ), //i
    .io_inputB               (pes_9_6_io_outputB[7:0]     ), //i
    .io_inputC               (pes_9_7_io_outputC[25:0]    ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_10_6), //i
    .io_resetPartialC        (io_resetPartialC_10_6       ), //i
    .io_outputA              (pes_10_6_io_outputA[7:0]    ), //o
    .io_outputB              (pes_10_6_io_outputB[7:0]    ), //o
    .io_outputC              (pes_10_6_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_10_7 (
    .io_inputA               (pes_10_6_io_outputA[7:0]    ), //i
    .io_inputB               (pes_9_7_io_outputB[7:0]     ), //i
    .io_inputC               (pes_9_8_io_outputC[25:0]    ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_10_7), //i
    .io_resetPartialC        (io_resetPartialC_10_7       ), //i
    .io_outputA              (pes_10_7_io_outputA[7:0]    ), //o
    .io_outputB              (pes_10_7_io_outputB[7:0]    ), //o
    .io_outputC              (pes_10_7_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_10_8 (
    .io_inputA               (pes_10_7_io_outputA[7:0]    ), //i
    .io_inputB               (pes_9_8_io_outputB[7:0]     ), //i
    .io_inputC               (pes_9_9_io_outputC[25:0]    ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_10_8), //i
    .io_resetPartialC        (io_resetPartialC_10_8       ), //i
    .io_outputA              (pes_10_8_io_outputA[7:0]    ), //o
    .io_outputB              (pes_10_8_io_outputB[7:0]    ), //o
    .io_outputC              (pes_10_8_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_10_9 (
    .io_inputA               (pes_10_8_io_outputA[7:0]    ), //i
    .io_inputB               (pes_9_9_io_outputB[7:0]     ), //i
    .io_inputC               (pes_9_10_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_10_9), //i
    .io_resetPartialC        (io_resetPartialC_10_9       ), //i
    .io_outputA              (pes_10_9_io_outputA[7:0]    ), //o
    .io_outputB              (pes_10_9_io_outputB[7:0]    ), //o
    .io_outputC              (pes_10_9_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_10_10 (
    .io_inputA               (pes_10_9_io_outputA[7:0]     ), //i
    .io_inputB               (pes_9_10_io_outputB[7:0]     ), //i
    .io_inputC               (pes_9_11_io_outputC[25:0]    ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_10_10), //i
    .io_resetPartialC        (io_resetPartialC_10_10       ), //i
    .io_outputA              (pes_10_10_io_outputA[7:0]    ), //o
    .io_outputB              (pes_10_10_io_outputB[7:0]    ), //o
    .io_outputC              (pes_10_10_io_outputC[25:0]   ), //o
    .clk                     (clk                          ), //i
    .reset                   (reset                        )  //i
  );
  ProcessingElement_16 pes_10_11 (
    .io_inputA               (pes_10_10_io_outputA[7:0]    ), //i
    .io_inputB               (pes_9_11_io_outputB[7:0]     ), //i
    .io_inputC               (pes_9_12_io_outputC[25:0]    ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_10_11), //i
    .io_resetPartialC        (io_resetPartialC_10_11       ), //i
    .io_outputA              (pes_10_11_io_outputA[7:0]    ), //o
    .io_outputB              (pes_10_11_io_outputB[7:0]    ), //o
    .io_outputC              (pes_10_11_io_outputC[25:0]   ), //o
    .clk                     (clk                          ), //i
    .reset                   (reset                        )  //i
  );
  ProcessingElement_16 pes_10_12 (
    .io_inputA               (pes_10_11_io_outputA[7:0]    ), //i
    .io_inputB               (pes_9_12_io_outputB[7:0]     ), //i
    .io_inputC               (pes_9_13_io_outputC[25:0]    ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_10_12), //i
    .io_resetPartialC        (io_resetPartialC_10_12       ), //i
    .io_outputA              (pes_10_12_io_outputA[7:0]    ), //o
    .io_outputB              (pes_10_12_io_outputB[7:0]    ), //o
    .io_outputC              (pes_10_12_io_outputC[25:0]   ), //o
    .clk                     (clk                          ), //i
    .reset                   (reset                        )  //i
  );
  ProcessingElement_16 pes_10_13 (
    .io_inputA               (pes_10_12_io_outputA[7:0]    ), //i
    .io_inputB               (pes_9_13_io_outputB[7:0]     ), //i
    .io_inputC               (pes_9_14_io_outputC[25:0]    ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_10_13), //i
    .io_resetPartialC        (io_resetPartialC_10_13       ), //i
    .io_outputA              (pes_10_13_io_outputA[7:0]    ), //o
    .io_outputB              (pes_10_13_io_outputB[7:0]    ), //o
    .io_outputC              (pes_10_13_io_outputC[25:0]   ), //o
    .clk                     (clk                          ), //i
    .reset                   (reset                        )  //i
  );
  ProcessingElement_16 pes_10_14 (
    .io_inputA               (pes_10_13_io_outputA[7:0]    ), //i
    .io_inputB               (pes_9_14_io_outputB[7:0]     ), //i
    .io_inputC               (pes_9_15_io_outputC[25:0]    ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_10_14), //i
    .io_resetPartialC        (io_resetPartialC_10_14       ), //i
    .io_outputA              (pes_10_14_io_outputA[7:0]    ), //o
    .io_outputB              (pes_10_14_io_outputB[7:0]    ), //o
    .io_outputC              (pes_10_14_io_outputC[25:0]   ), //o
    .clk                     (clk                          ), //i
    .reset                   (reset                        )  //i
  );
  ProcessingElement_15 pes_10_15 (
    .io_inputA               (pes_10_14_io_outputA[7:0]    ), //i
    .io_inputB               (pes_9_15_io_outputB[7:0]     ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_10_15), //i
    .io_resetPartialC        (io_resetPartialC_10_15       ), //i
    .io_outputB              (pes_10_15_io_outputB[7:0]    ), //o
    .io_outputC              (pes_10_15_io_outputC[25:0]   ), //o
    .clk                     (clk                          ), //i
    .reset                   (reset                        )  //i
  );
  ProcessingElement_16 pes_11_0 (
    .io_inputA               (skewBuffer_io_output_11[7:0]), //i
    .io_inputB               (pes_10_0_io_outputB[7:0]    ), //i
    .io_inputC               (pes_10_1_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_11_0), //i
    .io_resetPartialC        (io_resetPartialC_11_0       ), //i
    .io_outputA              (pes_11_0_io_outputA[7:0]    ), //o
    .io_outputB              (pes_11_0_io_outputB[7:0]    ), //o
    .io_outputC              (pes_11_0_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_11_1 (
    .io_inputA               (pes_11_0_io_outputA[7:0]    ), //i
    .io_inputB               (pes_10_1_io_outputB[7:0]    ), //i
    .io_inputC               (pes_10_2_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_11_1), //i
    .io_resetPartialC        (io_resetPartialC_11_1       ), //i
    .io_outputA              (pes_11_1_io_outputA[7:0]    ), //o
    .io_outputB              (pes_11_1_io_outputB[7:0]    ), //o
    .io_outputC              (pes_11_1_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_11_2 (
    .io_inputA               (pes_11_1_io_outputA[7:0]    ), //i
    .io_inputB               (pes_10_2_io_outputB[7:0]    ), //i
    .io_inputC               (pes_10_3_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_11_2), //i
    .io_resetPartialC        (io_resetPartialC_11_2       ), //i
    .io_outputA              (pes_11_2_io_outputA[7:0]    ), //o
    .io_outputB              (pes_11_2_io_outputB[7:0]    ), //o
    .io_outputC              (pes_11_2_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_11_3 (
    .io_inputA               (pes_11_2_io_outputA[7:0]    ), //i
    .io_inputB               (pes_10_3_io_outputB[7:0]    ), //i
    .io_inputC               (pes_10_4_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_11_3), //i
    .io_resetPartialC        (io_resetPartialC_11_3       ), //i
    .io_outputA              (pes_11_3_io_outputA[7:0]    ), //o
    .io_outputB              (pes_11_3_io_outputB[7:0]    ), //o
    .io_outputC              (pes_11_3_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_11_4 (
    .io_inputA               (pes_11_3_io_outputA[7:0]    ), //i
    .io_inputB               (pes_10_4_io_outputB[7:0]    ), //i
    .io_inputC               (pes_10_5_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_11_4), //i
    .io_resetPartialC        (io_resetPartialC_11_4       ), //i
    .io_outputA              (pes_11_4_io_outputA[7:0]    ), //o
    .io_outputB              (pes_11_4_io_outputB[7:0]    ), //o
    .io_outputC              (pes_11_4_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_11_5 (
    .io_inputA               (pes_11_4_io_outputA[7:0]    ), //i
    .io_inputB               (pes_10_5_io_outputB[7:0]    ), //i
    .io_inputC               (pes_10_6_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_11_5), //i
    .io_resetPartialC        (io_resetPartialC_11_5       ), //i
    .io_outputA              (pes_11_5_io_outputA[7:0]    ), //o
    .io_outputB              (pes_11_5_io_outputB[7:0]    ), //o
    .io_outputC              (pes_11_5_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_11_6 (
    .io_inputA               (pes_11_5_io_outputA[7:0]    ), //i
    .io_inputB               (pes_10_6_io_outputB[7:0]    ), //i
    .io_inputC               (pes_10_7_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_11_6), //i
    .io_resetPartialC        (io_resetPartialC_11_6       ), //i
    .io_outputA              (pes_11_6_io_outputA[7:0]    ), //o
    .io_outputB              (pes_11_6_io_outputB[7:0]    ), //o
    .io_outputC              (pes_11_6_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_11_7 (
    .io_inputA               (pes_11_6_io_outputA[7:0]    ), //i
    .io_inputB               (pes_10_7_io_outputB[7:0]    ), //i
    .io_inputC               (pes_10_8_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_11_7), //i
    .io_resetPartialC        (io_resetPartialC_11_7       ), //i
    .io_outputA              (pes_11_7_io_outputA[7:0]    ), //o
    .io_outputB              (pes_11_7_io_outputB[7:0]    ), //o
    .io_outputC              (pes_11_7_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_11_8 (
    .io_inputA               (pes_11_7_io_outputA[7:0]    ), //i
    .io_inputB               (pes_10_8_io_outputB[7:0]    ), //i
    .io_inputC               (pes_10_9_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_11_8), //i
    .io_resetPartialC        (io_resetPartialC_11_8       ), //i
    .io_outputA              (pes_11_8_io_outputA[7:0]    ), //o
    .io_outputB              (pes_11_8_io_outputB[7:0]    ), //o
    .io_outputC              (pes_11_8_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_11_9 (
    .io_inputA               (pes_11_8_io_outputA[7:0]    ), //i
    .io_inputB               (pes_10_9_io_outputB[7:0]    ), //i
    .io_inputC               (pes_10_10_io_outputC[25:0]  ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_11_9), //i
    .io_resetPartialC        (io_resetPartialC_11_9       ), //i
    .io_outputA              (pes_11_9_io_outputA[7:0]    ), //o
    .io_outputB              (pes_11_9_io_outputB[7:0]    ), //o
    .io_outputC              (pes_11_9_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_11_10 (
    .io_inputA               (pes_11_9_io_outputA[7:0]     ), //i
    .io_inputB               (pes_10_10_io_outputB[7:0]    ), //i
    .io_inputC               (pes_10_11_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_11_10), //i
    .io_resetPartialC        (io_resetPartialC_11_10       ), //i
    .io_outputA              (pes_11_10_io_outputA[7:0]    ), //o
    .io_outputB              (pes_11_10_io_outputB[7:0]    ), //o
    .io_outputC              (pes_11_10_io_outputC[25:0]   ), //o
    .clk                     (clk                          ), //i
    .reset                   (reset                        )  //i
  );
  ProcessingElement_16 pes_11_11 (
    .io_inputA               (pes_11_10_io_outputA[7:0]    ), //i
    .io_inputB               (pes_10_11_io_outputB[7:0]    ), //i
    .io_inputC               (pes_10_12_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_11_11), //i
    .io_resetPartialC        (io_resetPartialC_11_11       ), //i
    .io_outputA              (pes_11_11_io_outputA[7:0]    ), //o
    .io_outputB              (pes_11_11_io_outputB[7:0]    ), //o
    .io_outputC              (pes_11_11_io_outputC[25:0]   ), //o
    .clk                     (clk                          ), //i
    .reset                   (reset                        )  //i
  );
  ProcessingElement_16 pes_11_12 (
    .io_inputA               (pes_11_11_io_outputA[7:0]    ), //i
    .io_inputB               (pes_10_12_io_outputB[7:0]    ), //i
    .io_inputC               (pes_10_13_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_11_12), //i
    .io_resetPartialC        (io_resetPartialC_11_12       ), //i
    .io_outputA              (pes_11_12_io_outputA[7:0]    ), //o
    .io_outputB              (pes_11_12_io_outputB[7:0]    ), //o
    .io_outputC              (pes_11_12_io_outputC[25:0]   ), //o
    .clk                     (clk                          ), //i
    .reset                   (reset                        )  //i
  );
  ProcessingElement_16 pes_11_13 (
    .io_inputA               (pes_11_12_io_outputA[7:0]    ), //i
    .io_inputB               (pes_10_13_io_outputB[7:0]    ), //i
    .io_inputC               (pes_10_14_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_11_13), //i
    .io_resetPartialC        (io_resetPartialC_11_13       ), //i
    .io_outputA              (pes_11_13_io_outputA[7:0]    ), //o
    .io_outputB              (pes_11_13_io_outputB[7:0]    ), //o
    .io_outputC              (pes_11_13_io_outputC[25:0]   ), //o
    .clk                     (clk                          ), //i
    .reset                   (reset                        )  //i
  );
  ProcessingElement_16 pes_11_14 (
    .io_inputA               (pes_11_13_io_outputA[7:0]    ), //i
    .io_inputB               (pes_10_14_io_outputB[7:0]    ), //i
    .io_inputC               (pes_10_15_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_11_14), //i
    .io_resetPartialC        (io_resetPartialC_11_14       ), //i
    .io_outputA              (pes_11_14_io_outputA[7:0]    ), //o
    .io_outputB              (pes_11_14_io_outputB[7:0]    ), //o
    .io_outputC              (pes_11_14_io_outputC[25:0]   ), //o
    .clk                     (clk                          ), //i
    .reset                   (reset                        )  //i
  );
  ProcessingElement_15 pes_11_15 (
    .io_inputA               (pes_11_14_io_outputA[7:0]    ), //i
    .io_inputB               (pes_10_15_io_outputB[7:0]    ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_11_15), //i
    .io_resetPartialC        (io_resetPartialC_11_15       ), //i
    .io_outputB              (pes_11_15_io_outputB[7:0]    ), //o
    .io_outputC              (pes_11_15_io_outputC[25:0]   ), //o
    .clk                     (clk                          ), //i
    .reset                   (reset                        )  //i
  );
  ProcessingElement_16 pes_12_0 (
    .io_inputA               (skewBuffer_io_output_12[7:0]), //i
    .io_inputB               (pes_11_0_io_outputB[7:0]    ), //i
    .io_inputC               (pes_11_1_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_12_0), //i
    .io_resetPartialC        (io_resetPartialC_12_0       ), //i
    .io_outputA              (pes_12_0_io_outputA[7:0]    ), //o
    .io_outputB              (pes_12_0_io_outputB[7:0]    ), //o
    .io_outputC              (pes_12_0_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_12_1 (
    .io_inputA               (pes_12_0_io_outputA[7:0]    ), //i
    .io_inputB               (pes_11_1_io_outputB[7:0]    ), //i
    .io_inputC               (pes_11_2_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_12_1), //i
    .io_resetPartialC        (io_resetPartialC_12_1       ), //i
    .io_outputA              (pes_12_1_io_outputA[7:0]    ), //o
    .io_outputB              (pes_12_1_io_outputB[7:0]    ), //o
    .io_outputC              (pes_12_1_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_12_2 (
    .io_inputA               (pes_12_1_io_outputA[7:0]    ), //i
    .io_inputB               (pes_11_2_io_outputB[7:0]    ), //i
    .io_inputC               (pes_11_3_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_12_2), //i
    .io_resetPartialC        (io_resetPartialC_12_2       ), //i
    .io_outputA              (pes_12_2_io_outputA[7:0]    ), //o
    .io_outputB              (pes_12_2_io_outputB[7:0]    ), //o
    .io_outputC              (pes_12_2_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_12_3 (
    .io_inputA               (pes_12_2_io_outputA[7:0]    ), //i
    .io_inputB               (pes_11_3_io_outputB[7:0]    ), //i
    .io_inputC               (pes_11_4_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_12_3), //i
    .io_resetPartialC        (io_resetPartialC_12_3       ), //i
    .io_outputA              (pes_12_3_io_outputA[7:0]    ), //o
    .io_outputB              (pes_12_3_io_outputB[7:0]    ), //o
    .io_outputC              (pes_12_3_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_12_4 (
    .io_inputA               (pes_12_3_io_outputA[7:0]    ), //i
    .io_inputB               (pes_11_4_io_outputB[7:0]    ), //i
    .io_inputC               (pes_11_5_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_12_4), //i
    .io_resetPartialC        (io_resetPartialC_12_4       ), //i
    .io_outputA              (pes_12_4_io_outputA[7:0]    ), //o
    .io_outputB              (pes_12_4_io_outputB[7:0]    ), //o
    .io_outputC              (pes_12_4_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_12_5 (
    .io_inputA               (pes_12_4_io_outputA[7:0]    ), //i
    .io_inputB               (pes_11_5_io_outputB[7:0]    ), //i
    .io_inputC               (pes_11_6_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_12_5), //i
    .io_resetPartialC        (io_resetPartialC_12_5       ), //i
    .io_outputA              (pes_12_5_io_outputA[7:0]    ), //o
    .io_outputB              (pes_12_5_io_outputB[7:0]    ), //o
    .io_outputC              (pes_12_5_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_12_6 (
    .io_inputA               (pes_12_5_io_outputA[7:0]    ), //i
    .io_inputB               (pes_11_6_io_outputB[7:0]    ), //i
    .io_inputC               (pes_11_7_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_12_6), //i
    .io_resetPartialC        (io_resetPartialC_12_6       ), //i
    .io_outputA              (pes_12_6_io_outputA[7:0]    ), //o
    .io_outputB              (pes_12_6_io_outputB[7:0]    ), //o
    .io_outputC              (pes_12_6_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_12_7 (
    .io_inputA               (pes_12_6_io_outputA[7:0]    ), //i
    .io_inputB               (pes_11_7_io_outputB[7:0]    ), //i
    .io_inputC               (pes_11_8_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_12_7), //i
    .io_resetPartialC        (io_resetPartialC_12_7       ), //i
    .io_outputA              (pes_12_7_io_outputA[7:0]    ), //o
    .io_outputB              (pes_12_7_io_outputB[7:0]    ), //o
    .io_outputC              (pes_12_7_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_12_8 (
    .io_inputA               (pes_12_7_io_outputA[7:0]    ), //i
    .io_inputB               (pes_11_8_io_outputB[7:0]    ), //i
    .io_inputC               (pes_11_9_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_12_8), //i
    .io_resetPartialC        (io_resetPartialC_12_8       ), //i
    .io_outputA              (pes_12_8_io_outputA[7:0]    ), //o
    .io_outputB              (pes_12_8_io_outputB[7:0]    ), //o
    .io_outputC              (pes_12_8_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_12_9 (
    .io_inputA               (pes_12_8_io_outputA[7:0]    ), //i
    .io_inputB               (pes_11_9_io_outputB[7:0]    ), //i
    .io_inputC               (pes_11_10_io_outputC[25:0]  ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_12_9), //i
    .io_resetPartialC        (io_resetPartialC_12_9       ), //i
    .io_outputA              (pes_12_9_io_outputA[7:0]    ), //o
    .io_outputB              (pes_12_9_io_outputB[7:0]    ), //o
    .io_outputC              (pes_12_9_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_12_10 (
    .io_inputA               (pes_12_9_io_outputA[7:0]     ), //i
    .io_inputB               (pes_11_10_io_outputB[7:0]    ), //i
    .io_inputC               (pes_11_11_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_12_10), //i
    .io_resetPartialC        (io_resetPartialC_12_10       ), //i
    .io_outputA              (pes_12_10_io_outputA[7:0]    ), //o
    .io_outputB              (pes_12_10_io_outputB[7:0]    ), //o
    .io_outputC              (pes_12_10_io_outputC[25:0]   ), //o
    .clk                     (clk                          ), //i
    .reset                   (reset                        )  //i
  );
  ProcessingElement_16 pes_12_11 (
    .io_inputA               (pes_12_10_io_outputA[7:0]    ), //i
    .io_inputB               (pes_11_11_io_outputB[7:0]    ), //i
    .io_inputC               (pes_11_12_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_12_11), //i
    .io_resetPartialC        (io_resetPartialC_12_11       ), //i
    .io_outputA              (pes_12_11_io_outputA[7:0]    ), //o
    .io_outputB              (pes_12_11_io_outputB[7:0]    ), //o
    .io_outputC              (pes_12_11_io_outputC[25:0]   ), //o
    .clk                     (clk                          ), //i
    .reset                   (reset                        )  //i
  );
  ProcessingElement_16 pes_12_12 (
    .io_inputA               (pes_12_11_io_outputA[7:0]    ), //i
    .io_inputB               (pes_11_12_io_outputB[7:0]    ), //i
    .io_inputC               (pes_11_13_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_12_12), //i
    .io_resetPartialC        (io_resetPartialC_12_12       ), //i
    .io_outputA              (pes_12_12_io_outputA[7:0]    ), //o
    .io_outputB              (pes_12_12_io_outputB[7:0]    ), //o
    .io_outputC              (pes_12_12_io_outputC[25:0]   ), //o
    .clk                     (clk                          ), //i
    .reset                   (reset                        )  //i
  );
  ProcessingElement_16 pes_12_13 (
    .io_inputA               (pes_12_12_io_outputA[7:0]    ), //i
    .io_inputB               (pes_11_13_io_outputB[7:0]    ), //i
    .io_inputC               (pes_11_14_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_12_13), //i
    .io_resetPartialC        (io_resetPartialC_12_13       ), //i
    .io_outputA              (pes_12_13_io_outputA[7:0]    ), //o
    .io_outputB              (pes_12_13_io_outputB[7:0]    ), //o
    .io_outputC              (pes_12_13_io_outputC[25:0]   ), //o
    .clk                     (clk                          ), //i
    .reset                   (reset                        )  //i
  );
  ProcessingElement_16 pes_12_14 (
    .io_inputA               (pes_12_13_io_outputA[7:0]    ), //i
    .io_inputB               (pes_11_14_io_outputB[7:0]    ), //i
    .io_inputC               (pes_11_15_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_12_14), //i
    .io_resetPartialC        (io_resetPartialC_12_14       ), //i
    .io_outputA              (pes_12_14_io_outputA[7:0]    ), //o
    .io_outputB              (pes_12_14_io_outputB[7:0]    ), //o
    .io_outputC              (pes_12_14_io_outputC[25:0]   ), //o
    .clk                     (clk                          ), //i
    .reset                   (reset                        )  //i
  );
  ProcessingElement_15 pes_12_15 (
    .io_inputA               (pes_12_14_io_outputA[7:0]    ), //i
    .io_inputB               (pes_11_15_io_outputB[7:0]    ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_12_15), //i
    .io_resetPartialC        (io_resetPartialC_12_15       ), //i
    .io_outputB              (pes_12_15_io_outputB[7:0]    ), //o
    .io_outputC              (pes_12_15_io_outputC[25:0]   ), //o
    .clk                     (clk                          ), //i
    .reset                   (reset                        )  //i
  );
  ProcessingElement_16 pes_13_0 (
    .io_inputA               (skewBuffer_io_output_13[7:0]), //i
    .io_inputB               (pes_12_0_io_outputB[7:0]    ), //i
    .io_inputC               (pes_12_1_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_13_0), //i
    .io_resetPartialC        (io_resetPartialC_13_0       ), //i
    .io_outputA              (pes_13_0_io_outputA[7:0]    ), //o
    .io_outputB              (pes_13_0_io_outputB[7:0]    ), //o
    .io_outputC              (pes_13_0_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_13_1 (
    .io_inputA               (pes_13_0_io_outputA[7:0]    ), //i
    .io_inputB               (pes_12_1_io_outputB[7:0]    ), //i
    .io_inputC               (pes_12_2_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_13_1), //i
    .io_resetPartialC        (io_resetPartialC_13_1       ), //i
    .io_outputA              (pes_13_1_io_outputA[7:0]    ), //o
    .io_outputB              (pes_13_1_io_outputB[7:0]    ), //o
    .io_outputC              (pes_13_1_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_13_2 (
    .io_inputA               (pes_13_1_io_outputA[7:0]    ), //i
    .io_inputB               (pes_12_2_io_outputB[7:0]    ), //i
    .io_inputC               (pes_12_3_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_13_2), //i
    .io_resetPartialC        (io_resetPartialC_13_2       ), //i
    .io_outputA              (pes_13_2_io_outputA[7:0]    ), //o
    .io_outputB              (pes_13_2_io_outputB[7:0]    ), //o
    .io_outputC              (pes_13_2_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_13_3 (
    .io_inputA               (pes_13_2_io_outputA[7:0]    ), //i
    .io_inputB               (pes_12_3_io_outputB[7:0]    ), //i
    .io_inputC               (pes_12_4_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_13_3), //i
    .io_resetPartialC        (io_resetPartialC_13_3       ), //i
    .io_outputA              (pes_13_3_io_outputA[7:0]    ), //o
    .io_outputB              (pes_13_3_io_outputB[7:0]    ), //o
    .io_outputC              (pes_13_3_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_13_4 (
    .io_inputA               (pes_13_3_io_outputA[7:0]    ), //i
    .io_inputB               (pes_12_4_io_outputB[7:0]    ), //i
    .io_inputC               (pes_12_5_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_13_4), //i
    .io_resetPartialC        (io_resetPartialC_13_4       ), //i
    .io_outputA              (pes_13_4_io_outputA[7:0]    ), //o
    .io_outputB              (pes_13_4_io_outputB[7:0]    ), //o
    .io_outputC              (pes_13_4_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_13_5 (
    .io_inputA               (pes_13_4_io_outputA[7:0]    ), //i
    .io_inputB               (pes_12_5_io_outputB[7:0]    ), //i
    .io_inputC               (pes_12_6_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_13_5), //i
    .io_resetPartialC        (io_resetPartialC_13_5       ), //i
    .io_outputA              (pes_13_5_io_outputA[7:0]    ), //o
    .io_outputB              (pes_13_5_io_outputB[7:0]    ), //o
    .io_outputC              (pes_13_5_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_13_6 (
    .io_inputA               (pes_13_5_io_outputA[7:0]    ), //i
    .io_inputB               (pes_12_6_io_outputB[7:0]    ), //i
    .io_inputC               (pes_12_7_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_13_6), //i
    .io_resetPartialC        (io_resetPartialC_13_6       ), //i
    .io_outputA              (pes_13_6_io_outputA[7:0]    ), //o
    .io_outputB              (pes_13_6_io_outputB[7:0]    ), //o
    .io_outputC              (pes_13_6_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_13_7 (
    .io_inputA               (pes_13_6_io_outputA[7:0]    ), //i
    .io_inputB               (pes_12_7_io_outputB[7:0]    ), //i
    .io_inputC               (pes_12_8_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_13_7), //i
    .io_resetPartialC        (io_resetPartialC_13_7       ), //i
    .io_outputA              (pes_13_7_io_outputA[7:0]    ), //o
    .io_outputB              (pes_13_7_io_outputB[7:0]    ), //o
    .io_outputC              (pes_13_7_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_13_8 (
    .io_inputA               (pes_13_7_io_outputA[7:0]    ), //i
    .io_inputB               (pes_12_8_io_outputB[7:0]    ), //i
    .io_inputC               (pes_12_9_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_13_8), //i
    .io_resetPartialC        (io_resetPartialC_13_8       ), //i
    .io_outputA              (pes_13_8_io_outputA[7:0]    ), //o
    .io_outputB              (pes_13_8_io_outputB[7:0]    ), //o
    .io_outputC              (pes_13_8_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_13_9 (
    .io_inputA               (pes_13_8_io_outputA[7:0]    ), //i
    .io_inputB               (pes_12_9_io_outputB[7:0]    ), //i
    .io_inputC               (pes_12_10_io_outputC[25:0]  ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_13_9), //i
    .io_resetPartialC        (io_resetPartialC_13_9       ), //i
    .io_outputA              (pes_13_9_io_outputA[7:0]    ), //o
    .io_outputB              (pes_13_9_io_outputB[7:0]    ), //o
    .io_outputC              (pes_13_9_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_13_10 (
    .io_inputA               (pes_13_9_io_outputA[7:0]     ), //i
    .io_inputB               (pes_12_10_io_outputB[7:0]    ), //i
    .io_inputC               (pes_12_11_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_13_10), //i
    .io_resetPartialC        (io_resetPartialC_13_10       ), //i
    .io_outputA              (pes_13_10_io_outputA[7:0]    ), //o
    .io_outputB              (pes_13_10_io_outputB[7:0]    ), //o
    .io_outputC              (pes_13_10_io_outputC[25:0]   ), //o
    .clk                     (clk                          ), //i
    .reset                   (reset                        )  //i
  );
  ProcessingElement_16 pes_13_11 (
    .io_inputA               (pes_13_10_io_outputA[7:0]    ), //i
    .io_inputB               (pes_12_11_io_outputB[7:0]    ), //i
    .io_inputC               (pes_12_12_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_13_11), //i
    .io_resetPartialC        (io_resetPartialC_13_11       ), //i
    .io_outputA              (pes_13_11_io_outputA[7:0]    ), //o
    .io_outputB              (pes_13_11_io_outputB[7:0]    ), //o
    .io_outputC              (pes_13_11_io_outputC[25:0]   ), //o
    .clk                     (clk                          ), //i
    .reset                   (reset                        )  //i
  );
  ProcessingElement_16 pes_13_12 (
    .io_inputA               (pes_13_11_io_outputA[7:0]    ), //i
    .io_inputB               (pes_12_12_io_outputB[7:0]    ), //i
    .io_inputC               (pes_12_13_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_13_12), //i
    .io_resetPartialC        (io_resetPartialC_13_12       ), //i
    .io_outputA              (pes_13_12_io_outputA[7:0]    ), //o
    .io_outputB              (pes_13_12_io_outputB[7:0]    ), //o
    .io_outputC              (pes_13_12_io_outputC[25:0]   ), //o
    .clk                     (clk                          ), //i
    .reset                   (reset                        )  //i
  );
  ProcessingElement_16 pes_13_13 (
    .io_inputA               (pes_13_12_io_outputA[7:0]    ), //i
    .io_inputB               (pes_12_13_io_outputB[7:0]    ), //i
    .io_inputC               (pes_12_14_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_13_13), //i
    .io_resetPartialC        (io_resetPartialC_13_13       ), //i
    .io_outputA              (pes_13_13_io_outputA[7:0]    ), //o
    .io_outputB              (pes_13_13_io_outputB[7:0]    ), //o
    .io_outputC              (pes_13_13_io_outputC[25:0]   ), //o
    .clk                     (clk                          ), //i
    .reset                   (reset                        )  //i
  );
  ProcessingElement_16 pes_13_14 (
    .io_inputA               (pes_13_13_io_outputA[7:0]    ), //i
    .io_inputB               (pes_12_14_io_outputB[7:0]    ), //i
    .io_inputC               (pes_12_15_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_13_14), //i
    .io_resetPartialC        (io_resetPartialC_13_14       ), //i
    .io_outputA              (pes_13_14_io_outputA[7:0]    ), //o
    .io_outputB              (pes_13_14_io_outputB[7:0]    ), //o
    .io_outputC              (pes_13_14_io_outputC[25:0]   ), //o
    .clk                     (clk                          ), //i
    .reset                   (reset                        )  //i
  );
  ProcessingElement_15 pes_13_15 (
    .io_inputA               (pes_13_14_io_outputA[7:0]    ), //i
    .io_inputB               (pes_12_15_io_outputB[7:0]    ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_13_15), //i
    .io_resetPartialC        (io_resetPartialC_13_15       ), //i
    .io_outputB              (pes_13_15_io_outputB[7:0]    ), //o
    .io_outputC              (pes_13_15_io_outputC[25:0]   ), //o
    .clk                     (clk                          ), //i
    .reset                   (reset                        )  //i
  );
  ProcessingElement_16 pes_14_0 (
    .io_inputA               (skewBuffer_io_output_14[7:0]), //i
    .io_inputB               (pes_13_0_io_outputB[7:0]    ), //i
    .io_inputC               (pes_13_1_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_14_0), //i
    .io_resetPartialC        (io_resetPartialC_14_0       ), //i
    .io_outputA              (pes_14_0_io_outputA[7:0]    ), //o
    .io_outputB              (pes_14_0_io_outputB[7:0]    ), //o
    .io_outputC              (pes_14_0_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_14_1 (
    .io_inputA               (pes_14_0_io_outputA[7:0]    ), //i
    .io_inputB               (pes_13_1_io_outputB[7:0]    ), //i
    .io_inputC               (pes_13_2_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_14_1), //i
    .io_resetPartialC        (io_resetPartialC_14_1       ), //i
    .io_outputA              (pes_14_1_io_outputA[7:0]    ), //o
    .io_outputB              (pes_14_1_io_outputB[7:0]    ), //o
    .io_outputC              (pes_14_1_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_14_2 (
    .io_inputA               (pes_14_1_io_outputA[7:0]    ), //i
    .io_inputB               (pes_13_2_io_outputB[7:0]    ), //i
    .io_inputC               (pes_13_3_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_14_2), //i
    .io_resetPartialC        (io_resetPartialC_14_2       ), //i
    .io_outputA              (pes_14_2_io_outputA[7:0]    ), //o
    .io_outputB              (pes_14_2_io_outputB[7:0]    ), //o
    .io_outputC              (pes_14_2_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_14_3 (
    .io_inputA               (pes_14_2_io_outputA[7:0]    ), //i
    .io_inputB               (pes_13_3_io_outputB[7:0]    ), //i
    .io_inputC               (pes_13_4_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_14_3), //i
    .io_resetPartialC        (io_resetPartialC_14_3       ), //i
    .io_outputA              (pes_14_3_io_outputA[7:0]    ), //o
    .io_outputB              (pes_14_3_io_outputB[7:0]    ), //o
    .io_outputC              (pes_14_3_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_14_4 (
    .io_inputA               (pes_14_3_io_outputA[7:0]    ), //i
    .io_inputB               (pes_13_4_io_outputB[7:0]    ), //i
    .io_inputC               (pes_13_5_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_14_4), //i
    .io_resetPartialC        (io_resetPartialC_14_4       ), //i
    .io_outputA              (pes_14_4_io_outputA[7:0]    ), //o
    .io_outputB              (pes_14_4_io_outputB[7:0]    ), //o
    .io_outputC              (pes_14_4_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_14_5 (
    .io_inputA               (pes_14_4_io_outputA[7:0]    ), //i
    .io_inputB               (pes_13_5_io_outputB[7:0]    ), //i
    .io_inputC               (pes_13_6_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_14_5), //i
    .io_resetPartialC        (io_resetPartialC_14_5       ), //i
    .io_outputA              (pes_14_5_io_outputA[7:0]    ), //o
    .io_outputB              (pes_14_5_io_outputB[7:0]    ), //o
    .io_outputC              (pes_14_5_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_14_6 (
    .io_inputA               (pes_14_5_io_outputA[7:0]    ), //i
    .io_inputB               (pes_13_6_io_outputB[7:0]    ), //i
    .io_inputC               (pes_13_7_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_14_6), //i
    .io_resetPartialC        (io_resetPartialC_14_6       ), //i
    .io_outputA              (pes_14_6_io_outputA[7:0]    ), //o
    .io_outputB              (pes_14_6_io_outputB[7:0]    ), //o
    .io_outputC              (pes_14_6_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_14_7 (
    .io_inputA               (pes_14_6_io_outputA[7:0]    ), //i
    .io_inputB               (pes_13_7_io_outputB[7:0]    ), //i
    .io_inputC               (pes_13_8_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_14_7), //i
    .io_resetPartialC        (io_resetPartialC_14_7       ), //i
    .io_outputA              (pes_14_7_io_outputA[7:0]    ), //o
    .io_outputB              (pes_14_7_io_outputB[7:0]    ), //o
    .io_outputC              (pes_14_7_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_14_8 (
    .io_inputA               (pes_14_7_io_outputA[7:0]    ), //i
    .io_inputB               (pes_13_8_io_outputB[7:0]    ), //i
    .io_inputC               (pes_13_9_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_14_8), //i
    .io_resetPartialC        (io_resetPartialC_14_8       ), //i
    .io_outputA              (pes_14_8_io_outputA[7:0]    ), //o
    .io_outputB              (pes_14_8_io_outputB[7:0]    ), //o
    .io_outputC              (pes_14_8_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_14_9 (
    .io_inputA               (pes_14_8_io_outputA[7:0]    ), //i
    .io_inputB               (pes_13_9_io_outputB[7:0]    ), //i
    .io_inputC               (pes_13_10_io_outputC[25:0]  ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_14_9), //i
    .io_resetPartialC        (io_resetPartialC_14_9       ), //i
    .io_outputA              (pes_14_9_io_outputA[7:0]    ), //o
    .io_outputB              (pes_14_9_io_outputB[7:0]    ), //o
    .io_outputC              (pes_14_9_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_16 pes_14_10 (
    .io_inputA               (pes_14_9_io_outputA[7:0]     ), //i
    .io_inputB               (pes_13_10_io_outputB[7:0]    ), //i
    .io_inputC               (pes_13_11_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_14_10), //i
    .io_resetPartialC        (io_resetPartialC_14_10       ), //i
    .io_outputA              (pes_14_10_io_outputA[7:0]    ), //o
    .io_outputB              (pes_14_10_io_outputB[7:0]    ), //o
    .io_outputC              (pes_14_10_io_outputC[25:0]   ), //o
    .clk                     (clk                          ), //i
    .reset                   (reset                        )  //i
  );
  ProcessingElement_16 pes_14_11 (
    .io_inputA               (pes_14_10_io_outputA[7:0]    ), //i
    .io_inputB               (pes_13_11_io_outputB[7:0]    ), //i
    .io_inputC               (pes_13_12_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_14_11), //i
    .io_resetPartialC        (io_resetPartialC_14_11       ), //i
    .io_outputA              (pes_14_11_io_outputA[7:0]    ), //o
    .io_outputB              (pes_14_11_io_outputB[7:0]    ), //o
    .io_outputC              (pes_14_11_io_outputC[25:0]   ), //o
    .clk                     (clk                          ), //i
    .reset                   (reset                        )  //i
  );
  ProcessingElement_16 pes_14_12 (
    .io_inputA               (pes_14_11_io_outputA[7:0]    ), //i
    .io_inputB               (pes_13_12_io_outputB[7:0]    ), //i
    .io_inputC               (pes_13_13_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_14_12), //i
    .io_resetPartialC        (io_resetPartialC_14_12       ), //i
    .io_outputA              (pes_14_12_io_outputA[7:0]    ), //o
    .io_outputB              (pes_14_12_io_outputB[7:0]    ), //o
    .io_outputC              (pes_14_12_io_outputC[25:0]   ), //o
    .clk                     (clk                          ), //i
    .reset                   (reset                        )  //i
  );
  ProcessingElement_16 pes_14_13 (
    .io_inputA               (pes_14_12_io_outputA[7:0]    ), //i
    .io_inputB               (pes_13_13_io_outputB[7:0]    ), //i
    .io_inputC               (pes_13_14_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_14_13), //i
    .io_resetPartialC        (io_resetPartialC_14_13       ), //i
    .io_outputA              (pes_14_13_io_outputA[7:0]    ), //o
    .io_outputB              (pes_14_13_io_outputB[7:0]    ), //o
    .io_outputC              (pes_14_13_io_outputC[25:0]   ), //o
    .clk                     (clk                          ), //i
    .reset                   (reset                        )  //i
  );
  ProcessingElement_16 pes_14_14 (
    .io_inputA               (pes_14_13_io_outputA[7:0]    ), //i
    .io_inputB               (pes_13_14_io_outputB[7:0]    ), //i
    .io_inputC               (pes_13_15_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_14_14), //i
    .io_resetPartialC        (io_resetPartialC_14_14       ), //i
    .io_outputA              (pes_14_14_io_outputA[7:0]    ), //o
    .io_outputB              (pes_14_14_io_outputB[7:0]    ), //o
    .io_outputC              (pes_14_14_io_outputC[25:0]   ), //o
    .clk                     (clk                          ), //i
    .reset                   (reset                        )  //i
  );
  ProcessingElement_15 pes_14_15 (
    .io_inputA               (pes_14_14_io_outputA[7:0]    ), //i
    .io_inputB               (pes_13_15_io_outputB[7:0]    ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_14_15), //i
    .io_resetPartialC        (io_resetPartialC_14_15       ), //i
    .io_outputB              (pes_14_15_io_outputB[7:0]    ), //o
    .io_outputC              (pes_14_15_io_outputC[25:0]   ), //o
    .clk                     (clk                          ), //i
    .reset                   (reset                        )  //i
  );
  ProcessingElement_240 pes_15_0 (
    .io_inputA               (skewBuffer_io_output_15[7:0]), //i
    .io_inputB               (pes_14_0_io_outputB[7:0]    ), //i
    .io_inputC               (pes_14_1_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_15_0), //i
    .io_resetPartialC        (io_resetPartialC_15_0       ), //i
    .io_outputA              (pes_15_0_io_outputA[7:0]    ), //o
    .io_outputC              (pes_15_0_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_240 pes_15_1 (
    .io_inputA               (pes_15_0_io_outputA[7:0]    ), //i
    .io_inputB               (pes_14_1_io_outputB[7:0]    ), //i
    .io_inputC               (pes_14_2_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_15_1), //i
    .io_resetPartialC        (io_resetPartialC_15_1       ), //i
    .io_outputA              (pes_15_1_io_outputA[7:0]    ), //o
    .io_outputC              (pes_15_1_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_240 pes_15_2 (
    .io_inputA               (pes_15_1_io_outputA[7:0]    ), //i
    .io_inputB               (pes_14_2_io_outputB[7:0]    ), //i
    .io_inputC               (pes_14_3_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_15_2), //i
    .io_resetPartialC        (io_resetPartialC_15_2       ), //i
    .io_outputA              (pes_15_2_io_outputA[7:0]    ), //o
    .io_outputC              (pes_15_2_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_240 pes_15_3 (
    .io_inputA               (pes_15_2_io_outputA[7:0]    ), //i
    .io_inputB               (pes_14_3_io_outputB[7:0]    ), //i
    .io_inputC               (pes_14_4_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_15_3), //i
    .io_resetPartialC        (io_resetPartialC_15_3       ), //i
    .io_outputA              (pes_15_3_io_outputA[7:0]    ), //o
    .io_outputC              (pes_15_3_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_240 pes_15_4 (
    .io_inputA               (pes_15_3_io_outputA[7:0]    ), //i
    .io_inputB               (pes_14_4_io_outputB[7:0]    ), //i
    .io_inputC               (pes_14_5_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_15_4), //i
    .io_resetPartialC        (io_resetPartialC_15_4       ), //i
    .io_outputA              (pes_15_4_io_outputA[7:0]    ), //o
    .io_outputC              (pes_15_4_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_240 pes_15_5 (
    .io_inputA               (pes_15_4_io_outputA[7:0]    ), //i
    .io_inputB               (pes_14_5_io_outputB[7:0]    ), //i
    .io_inputC               (pes_14_6_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_15_5), //i
    .io_resetPartialC        (io_resetPartialC_15_5       ), //i
    .io_outputA              (pes_15_5_io_outputA[7:0]    ), //o
    .io_outputC              (pes_15_5_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_240 pes_15_6 (
    .io_inputA               (pes_15_5_io_outputA[7:0]    ), //i
    .io_inputB               (pes_14_6_io_outputB[7:0]    ), //i
    .io_inputC               (pes_14_7_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_15_6), //i
    .io_resetPartialC        (io_resetPartialC_15_6       ), //i
    .io_outputA              (pes_15_6_io_outputA[7:0]    ), //o
    .io_outputC              (pes_15_6_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_240 pes_15_7 (
    .io_inputA               (pes_15_6_io_outputA[7:0]    ), //i
    .io_inputB               (pes_14_7_io_outputB[7:0]    ), //i
    .io_inputC               (pes_14_8_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_15_7), //i
    .io_resetPartialC        (io_resetPartialC_15_7       ), //i
    .io_outputA              (pes_15_7_io_outputA[7:0]    ), //o
    .io_outputC              (pes_15_7_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_240 pes_15_8 (
    .io_inputA               (pes_15_7_io_outputA[7:0]    ), //i
    .io_inputB               (pes_14_8_io_outputB[7:0]    ), //i
    .io_inputC               (pes_14_9_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_15_8), //i
    .io_resetPartialC        (io_resetPartialC_15_8       ), //i
    .io_outputA              (pes_15_8_io_outputA[7:0]    ), //o
    .io_outputC              (pes_15_8_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_240 pes_15_9 (
    .io_inputA               (pes_15_8_io_outputA[7:0]    ), //i
    .io_inputB               (pes_14_9_io_outputB[7:0]    ), //i
    .io_inputC               (pes_14_10_io_outputC[25:0]  ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_15_9), //i
    .io_resetPartialC        (io_resetPartialC_15_9       ), //i
    .io_outputA              (pes_15_9_io_outputA[7:0]    ), //o
    .io_outputC              (pes_15_9_io_outputC[25:0]   ), //o
    .clk                     (clk                         ), //i
    .reset                   (reset                       )  //i
  );
  ProcessingElement_240 pes_15_10 (
    .io_inputA               (pes_15_9_io_outputA[7:0]     ), //i
    .io_inputB               (pes_14_10_io_outputB[7:0]    ), //i
    .io_inputC               (pes_14_11_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_15_10), //i
    .io_resetPartialC        (io_resetPartialC_15_10       ), //i
    .io_outputA              (pes_15_10_io_outputA[7:0]    ), //o
    .io_outputC              (pes_15_10_io_outputC[25:0]   ), //o
    .clk                     (clk                          ), //i
    .reset                   (reset                        )  //i
  );
  ProcessingElement_240 pes_15_11 (
    .io_inputA               (pes_15_10_io_outputA[7:0]    ), //i
    .io_inputB               (pes_14_11_io_outputB[7:0]    ), //i
    .io_inputC               (pes_14_12_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_15_11), //i
    .io_resetPartialC        (io_resetPartialC_15_11       ), //i
    .io_outputA              (pes_15_11_io_outputA[7:0]    ), //o
    .io_outputC              (pes_15_11_io_outputC[25:0]   ), //o
    .clk                     (clk                          ), //i
    .reset                   (reset                        )  //i
  );
  ProcessingElement_240 pes_15_12 (
    .io_inputA               (pes_15_11_io_outputA[7:0]    ), //i
    .io_inputB               (pes_14_12_io_outputB[7:0]    ), //i
    .io_inputC               (pes_14_13_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_15_12), //i
    .io_resetPartialC        (io_resetPartialC_15_12       ), //i
    .io_outputA              (pes_15_12_io_outputA[7:0]    ), //o
    .io_outputC              (pes_15_12_io_outputC[25:0]   ), //o
    .clk                     (clk                          ), //i
    .reset                   (reset                        )  //i
  );
  ProcessingElement_240 pes_15_13 (
    .io_inputA               (pes_15_12_io_outputA[7:0]    ), //i
    .io_inputB               (pes_14_13_io_outputB[7:0]    ), //i
    .io_inputC               (pes_14_14_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_15_13), //i
    .io_resetPartialC        (io_resetPartialC_15_13       ), //i
    .io_outputA              (pes_15_13_io_outputA[7:0]    ), //o
    .io_outputC              (pes_15_13_io_outputC[25:0]   ), //o
    .clk                     (clk                          ), //i
    .reset                   (reset                        )  //i
  );
  ProcessingElement_240 pes_15_14 (
    .io_inputA               (pes_15_13_io_outputA[7:0]    ), //i
    .io_inputB               (pes_14_14_io_outputB[7:0]    ), //i
    .io_inputC               (pes_14_15_io_outputC[25:0]   ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_15_14), //i
    .io_resetPartialC        (io_resetPartialC_15_14       ), //i
    .io_outputA              (pes_15_14_io_outputA[7:0]    ), //o
    .io_outputC              (pes_15_14_io_outputC[25:0]   ), //o
    .clk                     (clk                          ), //i
    .reset                   (reset                        )  //i
  );
  ProcessingElement_255 pes_15_15 (
    .io_inputA               (pes_15_14_io_outputA[7:0]    ), //i
    .io_inputB               (pes_14_15_io_outputB[7:0]    ), //i
    .io_outputCaptureEnableC (io_outputCaptureEnableC_15_15), //i
    .io_resetPartialC        (io_resetPartialC_15_15       ), //i
    .io_outputC              (pes_15_15_io_outputC[25:0]   ), //o
    .clk                     (clk                          ), //i
    .reset                   (reset                        )  //i
  );
  TypeA_SkewBuffer skewBuffer (
    .io_input_0   (io_inputA_0[7:0]            ), //i
    .io_input_1   (io_inputA_1[7:0]            ), //i
    .io_input_2   (io_inputA_2[7:0]            ), //i
    .io_input_3   (io_inputA_3[7:0]            ), //i
    .io_input_4   (io_inputA_4[7:0]            ), //i
    .io_input_5   (io_inputA_5[7:0]            ), //i
    .io_input_6   (io_inputA_6[7:0]            ), //i
    .io_input_7   (io_inputA_7[7:0]            ), //i
    .io_input_8   (io_inputA_8[7:0]            ), //i
    .io_input_9   (io_inputA_9[7:0]            ), //i
    .io_input_10  (io_inputA_10[7:0]           ), //i
    .io_input_11  (io_inputA_11[7:0]           ), //i
    .io_input_12  (io_inputA_12[7:0]           ), //i
    .io_input_13  (io_inputA_13[7:0]           ), //i
    .io_input_14  (io_inputA_14[7:0]           ), //i
    .io_input_15  (io_inputA_15[7:0]           ), //i
    .io_output_0  (skewBuffer_io_output_0[7:0] ), //o
    .io_output_1  (skewBuffer_io_output_1[7:0] ), //o
    .io_output_2  (skewBuffer_io_output_2[7:0] ), //o
    .io_output_3  (skewBuffer_io_output_3[7:0] ), //o
    .io_output_4  (skewBuffer_io_output_4[7:0] ), //o
    .io_output_5  (skewBuffer_io_output_5[7:0] ), //o
    .io_output_6  (skewBuffer_io_output_6[7:0] ), //o
    .io_output_7  (skewBuffer_io_output_7[7:0] ), //o
    .io_output_8  (skewBuffer_io_output_8[7:0] ), //o
    .io_output_9  (skewBuffer_io_output_9[7:0] ), //o
    .io_output_10 (skewBuffer_io_output_10[7:0]), //o
    .io_output_11 (skewBuffer_io_output_11[7:0]), //o
    .io_output_12 (skewBuffer_io_output_12[7:0]), //o
    .io_output_13 (skewBuffer_io_output_13[7:0]), //o
    .io_output_14 (skewBuffer_io_output_14[7:0]), //o
    .io_output_15 (skewBuffer_io_output_15[7:0]), //o
    .clk          (clk                         ), //i
    .reset        (reset                       )  //i
  );
  TypeB_SkewBuffer skewBuffer_1 (
    .io_input_0   (io_inputB_0[7:0]              ), //i
    .io_input_1   (io_inputB_1[7:0]              ), //i
    .io_input_2   (io_inputB_2[7:0]              ), //i
    .io_input_3   (io_inputB_3[7:0]              ), //i
    .io_input_4   (io_inputB_4[7:0]              ), //i
    .io_input_5   (io_inputB_5[7:0]              ), //i
    .io_input_6   (io_inputB_6[7:0]              ), //i
    .io_input_7   (io_inputB_7[7:0]              ), //i
    .io_input_8   (io_inputB_8[7:0]              ), //i
    .io_input_9   (io_inputB_9[7:0]              ), //i
    .io_input_10  (io_inputB_10[7:0]             ), //i
    .io_input_11  (io_inputB_11[7:0]             ), //i
    .io_input_12  (io_inputB_12[7:0]             ), //i
    .io_input_13  (io_inputB_13[7:0]             ), //i
    .io_input_14  (io_inputB_14[7:0]             ), //i
    .io_input_15  (io_inputB_15[7:0]             ), //i
    .io_output_0  (skewBuffer_1_io_output_0[7:0] ), //o
    .io_output_1  (skewBuffer_1_io_output_1[7:0] ), //o
    .io_output_2  (skewBuffer_1_io_output_2[7:0] ), //o
    .io_output_3  (skewBuffer_1_io_output_3[7:0] ), //o
    .io_output_4  (skewBuffer_1_io_output_4[7:0] ), //o
    .io_output_5  (skewBuffer_1_io_output_5[7:0] ), //o
    .io_output_6  (skewBuffer_1_io_output_6[7:0] ), //o
    .io_output_7  (skewBuffer_1_io_output_7[7:0] ), //o
    .io_output_8  (skewBuffer_1_io_output_8[7:0] ), //o
    .io_output_9  (skewBuffer_1_io_output_9[7:0] ), //o
    .io_output_10 (skewBuffer_1_io_output_10[7:0]), //o
    .io_output_11 (skewBuffer_1_io_output_11[7:0]), //o
    .io_output_12 (skewBuffer_1_io_output_12[7:0]), //o
    .io_output_13 (skewBuffer_1_io_output_13[7:0]), //o
    .io_output_14 (skewBuffer_1_io_output_14[7:0]), //o
    .io_output_15 (skewBuffer_1_io_output_15[7:0]), //o
    .clk          (clk                           ), //i
    .reset        (reset                         )  //i
  );
  TypeC_DeskewBuffer deskewBufferReuseC (
    .io_input_0   (pes_0_0_io_outputC[25:0]             ), //i
    .io_input_1   (pes_1_0_io_outputC[25:0]             ), //i
    .io_input_2   (pes_2_0_io_outputC[25:0]             ), //i
    .io_input_3   (pes_3_0_io_outputC[25:0]             ), //i
    .io_input_4   (pes_4_0_io_outputC[25:0]             ), //i
    .io_input_5   (pes_5_0_io_outputC[25:0]             ), //i
    .io_input_6   (pes_6_0_io_outputC[25:0]             ), //i
    .io_input_7   (pes_7_0_io_outputC[25:0]             ), //i
    .io_input_8   (pes_8_0_io_outputC[25:0]             ), //i
    .io_input_9   (pes_9_0_io_outputC[25:0]             ), //i
    .io_input_10  (pes_10_0_io_outputC[25:0]            ), //i
    .io_input_11  (pes_11_0_io_outputC[25:0]            ), //i
    .io_input_12  (pes_12_0_io_outputC[25:0]            ), //i
    .io_input_13  (pes_13_0_io_outputC[25:0]            ), //i
    .io_input_14  (pes_14_0_io_outputC[25:0]            ), //i
    .io_input_15  (pes_15_0_io_outputC[25:0]            ), //i
    .io_input_16  (pes_15_1_io_outputC[25:0]            ), //i
    .io_input_17  (pes_15_2_io_outputC[25:0]            ), //i
    .io_input_18  (pes_15_3_io_outputC[25:0]            ), //i
    .io_input_19  (pes_15_4_io_outputC[25:0]            ), //i
    .io_input_20  (pes_15_5_io_outputC[25:0]            ), //i
    .io_input_21  (pes_15_6_io_outputC[25:0]            ), //i
    .io_input_22  (pes_15_7_io_outputC[25:0]            ), //i
    .io_input_23  (pes_15_8_io_outputC[25:0]            ), //i
    .io_input_24  (pes_15_9_io_outputC[25:0]            ), //i
    .io_input_25  (pes_15_10_io_outputC[25:0]           ), //i
    .io_input_26  (pes_15_11_io_outputC[25:0]           ), //i
    .io_input_27  (pes_15_12_io_outputC[25:0]           ), //i
    .io_input_28  (pes_15_13_io_outputC[25:0]           ), //i
    .io_input_29  (pes_15_14_io_outputC[25:0]           ), //i
    .io_input_30  (pes_15_15_io_outputC[25:0]           ), //i
    .io_output_0  (deskewBufferReuseC_io_output_0[25:0] ), //o
    .io_output_1  (deskewBufferReuseC_io_output_1[25:0] ), //o
    .io_output_2  (deskewBufferReuseC_io_output_2[25:0] ), //o
    .io_output_3  (deskewBufferReuseC_io_output_3[25:0] ), //o
    .io_output_4  (deskewBufferReuseC_io_output_4[25:0] ), //o
    .io_output_5  (deskewBufferReuseC_io_output_5[25:0] ), //o
    .io_output_6  (deskewBufferReuseC_io_output_6[25:0] ), //o
    .io_output_7  (deskewBufferReuseC_io_output_7[25:0] ), //o
    .io_output_8  (deskewBufferReuseC_io_output_8[25:0] ), //o
    .io_output_9  (deskewBufferReuseC_io_output_9[25:0] ), //o
    .io_output_10 (deskewBufferReuseC_io_output_10[25:0]), //o
    .io_output_11 (deskewBufferReuseC_io_output_11[25:0]), //o
    .io_output_12 (deskewBufferReuseC_io_output_12[25:0]), //o
    .io_output_13 (deskewBufferReuseC_io_output_13[25:0]), //o
    .io_output_14 (deskewBufferReuseC_io_output_14[25:0]), //o
    .io_output_15 (deskewBufferReuseC_io_output_15[25:0]), //o
    .io_output_16 (deskewBufferReuseC_io_output_16[25:0]), //o
    .io_output_17 (deskewBufferReuseC_io_output_17[25:0]), //o
    .io_output_18 (deskewBufferReuseC_io_output_18[25:0]), //o
    .io_output_19 (deskewBufferReuseC_io_output_19[25:0]), //o
    .io_output_20 (deskewBufferReuseC_io_output_20[25:0]), //o
    .io_output_21 (deskewBufferReuseC_io_output_21[25:0]), //o
    .io_output_22 (deskewBufferReuseC_io_output_22[25:0]), //o
    .io_output_23 (deskewBufferReuseC_io_output_23[25:0]), //o
    .io_output_24 (deskewBufferReuseC_io_output_24[25:0]), //o
    .io_output_25 (deskewBufferReuseC_io_output_25[25:0]), //o
    .io_output_26 (deskewBufferReuseC_io_output_26[25:0]), //o
    .io_output_27 (deskewBufferReuseC_io_output_27[25:0]), //o
    .io_output_28 (deskewBufferReuseC_io_output_28[25:0]), //o
    .io_output_29 (deskewBufferReuseC_io_output_29[25:0]), //o
    .io_output_30 (deskewBufferReuseC_io_output_30[25:0]), //o
    .clk          (clk                                  ), //i
    .reset        (reset                                )  //i
  );
  assign io_outputC_0 = deskewBufferReuseC_io_output_0;
  assign io_outputC_1 = deskewBufferReuseC_io_output_1;
  assign io_outputC_2 = deskewBufferReuseC_io_output_2;
  assign io_outputC_3 = deskewBufferReuseC_io_output_3;
  assign io_outputC_4 = deskewBufferReuseC_io_output_4;
  assign io_outputC_5 = deskewBufferReuseC_io_output_5;
  assign io_outputC_6 = deskewBufferReuseC_io_output_6;
  assign io_outputC_7 = deskewBufferReuseC_io_output_7;
  assign io_outputC_8 = deskewBufferReuseC_io_output_8;
  assign io_outputC_9 = deskewBufferReuseC_io_output_9;
  assign io_outputC_10 = deskewBufferReuseC_io_output_10;
  assign io_outputC_11 = deskewBufferReuseC_io_output_11;
  assign io_outputC_12 = deskewBufferReuseC_io_output_12;
  assign io_outputC_13 = deskewBufferReuseC_io_output_13;
  assign io_outputC_14 = deskewBufferReuseC_io_output_14;
  assign io_outputC_15 = deskewBufferReuseC_io_output_15;
  assign io_outputC_16 = deskewBufferReuseC_io_output_16;
  assign io_outputC_17 = deskewBufferReuseC_io_output_17;
  assign io_outputC_18 = deskewBufferReuseC_io_output_18;
  assign io_outputC_19 = deskewBufferReuseC_io_output_19;
  assign io_outputC_20 = deskewBufferReuseC_io_output_20;
  assign io_outputC_21 = deskewBufferReuseC_io_output_21;
  assign io_outputC_22 = deskewBufferReuseC_io_output_22;
  assign io_outputC_23 = deskewBufferReuseC_io_output_23;
  assign io_outputC_24 = deskewBufferReuseC_io_output_24;
  assign io_outputC_25 = deskewBufferReuseC_io_output_25;
  assign io_outputC_26 = deskewBufferReuseC_io_output_26;
  assign io_outputC_27 = deskewBufferReuseC_io_output_27;
  assign io_outputC_28 = deskewBufferReuseC_io_output_28;
  assign io_outputC_29 = deskewBufferReuseC_io_output_29;
  assign io_outputC_30 = deskewBufferReuseC_io_output_30;

endmodule

module TypeC_DeskewBuffer (
  input  wire [25:0]   io_input_0,
  input  wire [25:0]   io_input_1,
  input  wire [25:0]   io_input_2,
  input  wire [25:0]   io_input_3,
  input  wire [25:0]   io_input_4,
  input  wire [25:0]   io_input_5,
  input  wire [25:0]   io_input_6,
  input  wire [25:0]   io_input_7,
  input  wire [25:0]   io_input_8,
  input  wire [25:0]   io_input_9,
  input  wire [25:0]   io_input_10,
  input  wire [25:0]   io_input_11,
  input  wire [25:0]   io_input_12,
  input  wire [25:0]   io_input_13,
  input  wire [25:0]   io_input_14,
  input  wire [25:0]   io_input_15,
  input  wire [25:0]   io_input_16,
  input  wire [25:0]   io_input_17,
  input  wire [25:0]   io_input_18,
  input  wire [25:0]   io_input_19,
  input  wire [25:0]   io_input_20,
  input  wire [25:0]   io_input_21,
  input  wire [25:0]   io_input_22,
  input  wire [25:0]   io_input_23,
  input  wire [25:0]   io_input_24,
  input  wire [25:0]   io_input_25,
  input  wire [25:0]   io_input_26,
  input  wire [25:0]   io_input_27,
  input  wire [25:0]   io_input_28,
  input  wire [25:0]   io_input_29,
  input  wire [25:0]   io_input_30,
  output wire [25:0]   io_output_0,
  output wire [25:0]   io_output_1,
  output wire [25:0]   io_output_2,
  output wire [25:0]   io_output_3,
  output wire [25:0]   io_output_4,
  output wire [25:0]   io_output_5,
  output wire [25:0]   io_output_6,
  output wire [25:0]   io_output_7,
  output wire [25:0]   io_output_8,
  output wire [25:0]   io_output_9,
  output wire [25:0]   io_output_10,
  output wire [25:0]   io_output_11,
  output wire [25:0]   io_output_12,
  output wire [25:0]   io_output_13,
  output wire [25:0]   io_output_14,
  output wire [25:0]   io_output_15,
  output wire [25:0]   io_output_16,
  output wire [25:0]   io_output_17,
  output wire [25:0]   io_output_18,
  output wire [25:0]   io_output_19,
  output wire [25:0]   io_output_20,
  output wire [25:0]   io_output_21,
  output wire [25:0]   io_output_22,
  output wire [25:0]   io_output_23,
  output wire [25:0]   io_output_24,
  output wire [25:0]   io_output_25,
  output wire [25:0]   io_output_26,
  output wire [25:0]   io_output_27,
  output wire [25:0]   io_output_28,
  output wire [25:0]   io_output_29,
  output wire [25:0]   io_output_30,
  input  wire          clk,
  input  wire          reset
);

  reg        [25:0]   io_input_0_delay_1;
  reg        [25:0]   io_input_0_delay_2;
  reg        [25:0]   io_input_0_delay_3;
  reg        [25:0]   io_input_0_delay_4;
  reg        [25:0]   io_input_0_delay_5;
  reg        [25:0]   io_input_0_delay_6;
  reg        [25:0]   io_input_0_delay_7;
  reg        [25:0]   io_input_0_delay_8;
  reg        [25:0]   io_input_0_delay_9;
  reg        [25:0]   io_input_0_delay_10;
  reg        [25:0]   io_input_0_delay_11;
  reg        [25:0]   io_input_0_delay_12;
  reg        [25:0]   io_input_0_delay_13;
  reg        [25:0]   io_input_0_delay_14;
  reg        [25:0]   io_input_0_delay_15;
  reg        [25:0]   io_input_1_delay_1;
  reg        [25:0]   io_input_1_delay_2;
  reg        [25:0]   io_input_1_delay_3;
  reg        [25:0]   io_input_1_delay_4;
  reg        [25:0]   io_input_1_delay_5;
  reg        [25:0]   io_input_1_delay_6;
  reg        [25:0]   io_input_1_delay_7;
  reg        [25:0]   io_input_1_delay_8;
  reg        [25:0]   io_input_1_delay_9;
  reg        [25:0]   io_input_1_delay_10;
  reg        [25:0]   io_input_1_delay_11;
  reg        [25:0]   io_input_1_delay_12;
  reg        [25:0]   io_input_1_delay_13;
  reg        [25:0]   io_input_1_delay_14;
  reg        [25:0]   io_input_2_delay_1;
  reg        [25:0]   io_input_2_delay_2;
  reg        [25:0]   io_input_2_delay_3;
  reg        [25:0]   io_input_2_delay_4;
  reg        [25:0]   io_input_2_delay_5;
  reg        [25:0]   io_input_2_delay_6;
  reg        [25:0]   io_input_2_delay_7;
  reg        [25:0]   io_input_2_delay_8;
  reg        [25:0]   io_input_2_delay_9;
  reg        [25:0]   io_input_2_delay_10;
  reg        [25:0]   io_input_2_delay_11;
  reg        [25:0]   io_input_2_delay_12;
  reg        [25:0]   io_input_2_delay_13;
  reg        [25:0]   io_input_3_delay_1;
  reg        [25:0]   io_input_3_delay_2;
  reg        [25:0]   io_input_3_delay_3;
  reg        [25:0]   io_input_3_delay_4;
  reg        [25:0]   io_input_3_delay_5;
  reg        [25:0]   io_input_3_delay_6;
  reg        [25:0]   io_input_3_delay_7;
  reg        [25:0]   io_input_3_delay_8;
  reg        [25:0]   io_input_3_delay_9;
  reg        [25:0]   io_input_3_delay_10;
  reg        [25:0]   io_input_3_delay_11;
  reg        [25:0]   io_input_3_delay_12;
  reg        [25:0]   io_input_4_delay_1;
  reg        [25:0]   io_input_4_delay_2;
  reg        [25:0]   io_input_4_delay_3;
  reg        [25:0]   io_input_4_delay_4;
  reg        [25:0]   io_input_4_delay_5;
  reg        [25:0]   io_input_4_delay_6;
  reg        [25:0]   io_input_4_delay_7;
  reg        [25:0]   io_input_4_delay_8;
  reg        [25:0]   io_input_4_delay_9;
  reg        [25:0]   io_input_4_delay_10;
  reg        [25:0]   io_input_4_delay_11;
  reg        [25:0]   io_input_5_delay_1;
  reg        [25:0]   io_input_5_delay_2;
  reg        [25:0]   io_input_5_delay_3;
  reg        [25:0]   io_input_5_delay_4;
  reg        [25:0]   io_input_5_delay_5;
  reg        [25:0]   io_input_5_delay_6;
  reg        [25:0]   io_input_5_delay_7;
  reg        [25:0]   io_input_5_delay_8;
  reg        [25:0]   io_input_5_delay_9;
  reg        [25:0]   io_input_5_delay_10;
  reg        [25:0]   io_input_6_delay_1;
  reg        [25:0]   io_input_6_delay_2;
  reg        [25:0]   io_input_6_delay_3;
  reg        [25:0]   io_input_6_delay_4;
  reg        [25:0]   io_input_6_delay_5;
  reg        [25:0]   io_input_6_delay_6;
  reg        [25:0]   io_input_6_delay_7;
  reg        [25:0]   io_input_6_delay_8;
  reg        [25:0]   io_input_6_delay_9;
  reg        [25:0]   io_input_7_delay_1;
  reg        [25:0]   io_input_7_delay_2;
  reg        [25:0]   io_input_7_delay_3;
  reg        [25:0]   io_input_7_delay_4;
  reg        [25:0]   io_input_7_delay_5;
  reg        [25:0]   io_input_7_delay_6;
  reg        [25:0]   io_input_7_delay_7;
  reg        [25:0]   io_input_7_delay_8;
  reg        [25:0]   io_input_8_delay_1;
  reg        [25:0]   io_input_8_delay_2;
  reg        [25:0]   io_input_8_delay_3;
  reg        [25:0]   io_input_8_delay_4;
  reg        [25:0]   io_input_8_delay_5;
  reg        [25:0]   io_input_8_delay_6;
  reg        [25:0]   io_input_8_delay_7;
  reg        [25:0]   io_input_9_delay_1;
  reg        [25:0]   io_input_9_delay_2;
  reg        [25:0]   io_input_9_delay_3;
  reg        [25:0]   io_input_9_delay_4;
  reg        [25:0]   io_input_9_delay_5;
  reg        [25:0]   io_input_9_delay_6;
  reg        [25:0]   io_input_10_delay_1;
  reg        [25:0]   io_input_10_delay_2;
  reg        [25:0]   io_input_10_delay_3;
  reg        [25:0]   io_input_10_delay_4;
  reg        [25:0]   io_input_10_delay_5;
  reg        [25:0]   io_input_11_delay_1;
  reg        [25:0]   io_input_11_delay_2;
  reg        [25:0]   io_input_11_delay_3;
  reg        [25:0]   io_input_11_delay_4;
  reg        [25:0]   io_input_12_delay_1;
  reg        [25:0]   io_input_12_delay_2;
  reg        [25:0]   io_input_12_delay_3;
  reg        [25:0]   io_input_13_delay_1;
  reg        [25:0]   io_input_13_delay_2;
  reg        [25:0]   io_input_14_delay_1;

  assign io_output_0 = io_input_0_delay_15;
  assign io_output_1 = io_input_1_delay_14;
  assign io_output_2 = io_input_2_delay_13;
  assign io_output_3 = io_input_3_delay_12;
  assign io_output_4 = io_input_4_delay_11;
  assign io_output_5 = io_input_5_delay_10;
  assign io_output_6 = io_input_6_delay_9;
  assign io_output_7 = io_input_7_delay_8;
  assign io_output_8 = io_input_8_delay_7;
  assign io_output_9 = io_input_9_delay_6;
  assign io_output_10 = io_input_10_delay_5;
  assign io_output_11 = io_input_11_delay_4;
  assign io_output_12 = io_input_12_delay_3;
  assign io_output_13 = io_input_13_delay_2;
  assign io_output_14 = io_input_14_delay_1;
  assign io_output_15 = io_input_15;
  assign io_output_16 = io_input_16;
  assign io_output_17 = io_input_17;
  assign io_output_18 = io_input_18;
  assign io_output_19 = io_input_19;
  assign io_output_20 = io_input_20;
  assign io_output_21 = io_input_21;
  assign io_output_22 = io_input_22;
  assign io_output_23 = io_input_23;
  assign io_output_24 = io_input_24;
  assign io_output_25 = io_input_25;
  assign io_output_26 = io_input_26;
  assign io_output_27 = io_input_27;
  assign io_output_28 = io_input_28;
  assign io_output_29 = io_input_29;
  assign io_output_30 = io_input_30;
  always @(posedge clk) begin
    io_input_0_delay_1 <= io_input_0;
    io_input_0_delay_2 <= io_input_0_delay_1;
    io_input_0_delay_3 <= io_input_0_delay_2;
    io_input_0_delay_4 <= io_input_0_delay_3;
    io_input_0_delay_5 <= io_input_0_delay_4;
    io_input_0_delay_6 <= io_input_0_delay_5;
    io_input_0_delay_7 <= io_input_0_delay_6;
    io_input_0_delay_8 <= io_input_0_delay_7;
    io_input_0_delay_9 <= io_input_0_delay_8;
    io_input_0_delay_10 <= io_input_0_delay_9;
    io_input_0_delay_11 <= io_input_0_delay_10;
    io_input_0_delay_12 <= io_input_0_delay_11;
    io_input_0_delay_13 <= io_input_0_delay_12;
    io_input_0_delay_14 <= io_input_0_delay_13;
    io_input_0_delay_15 <= io_input_0_delay_14;
    io_input_1_delay_1 <= io_input_1;
    io_input_1_delay_2 <= io_input_1_delay_1;
    io_input_1_delay_3 <= io_input_1_delay_2;
    io_input_1_delay_4 <= io_input_1_delay_3;
    io_input_1_delay_5 <= io_input_1_delay_4;
    io_input_1_delay_6 <= io_input_1_delay_5;
    io_input_1_delay_7 <= io_input_1_delay_6;
    io_input_1_delay_8 <= io_input_1_delay_7;
    io_input_1_delay_9 <= io_input_1_delay_8;
    io_input_1_delay_10 <= io_input_1_delay_9;
    io_input_1_delay_11 <= io_input_1_delay_10;
    io_input_1_delay_12 <= io_input_1_delay_11;
    io_input_1_delay_13 <= io_input_1_delay_12;
    io_input_1_delay_14 <= io_input_1_delay_13;
    io_input_2_delay_1 <= io_input_2;
    io_input_2_delay_2 <= io_input_2_delay_1;
    io_input_2_delay_3 <= io_input_2_delay_2;
    io_input_2_delay_4 <= io_input_2_delay_3;
    io_input_2_delay_5 <= io_input_2_delay_4;
    io_input_2_delay_6 <= io_input_2_delay_5;
    io_input_2_delay_7 <= io_input_2_delay_6;
    io_input_2_delay_8 <= io_input_2_delay_7;
    io_input_2_delay_9 <= io_input_2_delay_8;
    io_input_2_delay_10 <= io_input_2_delay_9;
    io_input_2_delay_11 <= io_input_2_delay_10;
    io_input_2_delay_12 <= io_input_2_delay_11;
    io_input_2_delay_13 <= io_input_2_delay_12;
    io_input_3_delay_1 <= io_input_3;
    io_input_3_delay_2 <= io_input_3_delay_1;
    io_input_3_delay_3 <= io_input_3_delay_2;
    io_input_3_delay_4 <= io_input_3_delay_3;
    io_input_3_delay_5 <= io_input_3_delay_4;
    io_input_3_delay_6 <= io_input_3_delay_5;
    io_input_3_delay_7 <= io_input_3_delay_6;
    io_input_3_delay_8 <= io_input_3_delay_7;
    io_input_3_delay_9 <= io_input_3_delay_8;
    io_input_3_delay_10 <= io_input_3_delay_9;
    io_input_3_delay_11 <= io_input_3_delay_10;
    io_input_3_delay_12 <= io_input_3_delay_11;
    io_input_4_delay_1 <= io_input_4;
    io_input_4_delay_2 <= io_input_4_delay_1;
    io_input_4_delay_3 <= io_input_4_delay_2;
    io_input_4_delay_4 <= io_input_4_delay_3;
    io_input_4_delay_5 <= io_input_4_delay_4;
    io_input_4_delay_6 <= io_input_4_delay_5;
    io_input_4_delay_7 <= io_input_4_delay_6;
    io_input_4_delay_8 <= io_input_4_delay_7;
    io_input_4_delay_9 <= io_input_4_delay_8;
    io_input_4_delay_10 <= io_input_4_delay_9;
    io_input_4_delay_11 <= io_input_4_delay_10;
    io_input_5_delay_1 <= io_input_5;
    io_input_5_delay_2 <= io_input_5_delay_1;
    io_input_5_delay_3 <= io_input_5_delay_2;
    io_input_5_delay_4 <= io_input_5_delay_3;
    io_input_5_delay_5 <= io_input_5_delay_4;
    io_input_5_delay_6 <= io_input_5_delay_5;
    io_input_5_delay_7 <= io_input_5_delay_6;
    io_input_5_delay_8 <= io_input_5_delay_7;
    io_input_5_delay_9 <= io_input_5_delay_8;
    io_input_5_delay_10 <= io_input_5_delay_9;
    io_input_6_delay_1 <= io_input_6;
    io_input_6_delay_2 <= io_input_6_delay_1;
    io_input_6_delay_3 <= io_input_6_delay_2;
    io_input_6_delay_4 <= io_input_6_delay_3;
    io_input_6_delay_5 <= io_input_6_delay_4;
    io_input_6_delay_6 <= io_input_6_delay_5;
    io_input_6_delay_7 <= io_input_6_delay_6;
    io_input_6_delay_8 <= io_input_6_delay_7;
    io_input_6_delay_9 <= io_input_6_delay_8;
    io_input_7_delay_1 <= io_input_7;
    io_input_7_delay_2 <= io_input_7_delay_1;
    io_input_7_delay_3 <= io_input_7_delay_2;
    io_input_7_delay_4 <= io_input_7_delay_3;
    io_input_7_delay_5 <= io_input_7_delay_4;
    io_input_7_delay_6 <= io_input_7_delay_5;
    io_input_7_delay_7 <= io_input_7_delay_6;
    io_input_7_delay_8 <= io_input_7_delay_7;
    io_input_8_delay_1 <= io_input_8;
    io_input_8_delay_2 <= io_input_8_delay_1;
    io_input_8_delay_3 <= io_input_8_delay_2;
    io_input_8_delay_4 <= io_input_8_delay_3;
    io_input_8_delay_5 <= io_input_8_delay_4;
    io_input_8_delay_6 <= io_input_8_delay_5;
    io_input_8_delay_7 <= io_input_8_delay_6;
    io_input_9_delay_1 <= io_input_9;
    io_input_9_delay_2 <= io_input_9_delay_1;
    io_input_9_delay_3 <= io_input_9_delay_2;
    io_input_9_delay_4 <= io_input_9_delay_3;
    io_input_9_delay_5 <= io_input_9_delay_4;
    io_input_9_delay_6 <= io_input_9_delay_5;
    io_input_10_delay_1 <= io_input_10;
    io_input_10_delay_2 <= io_input_10_delay_1;
    io_input_10_delay_3 <= io_input_10_delay_2;
    io_input_10_delay_4 <= io_input_10_delay_3;
    io_input_10_delay_5 <= io_input_10_delay_4;
    io_input_11_delay_1 <= io_input_11;
    io_input_11_delay_2 <= io_input_11_delay_1;
    io_input_11_delay_3 <= io_input_11_delay_2;
    io_input_11_delay_4 <= io_input_11_delay_3;
    io_input_12_delay_1 <= io_input_12;
    io_input_12_delay_2 <= io_input_12_delay_1;
    io_input_12_delay_3 <= io_input_12_delay_2;
    io_input_13_delay_1 <= io_input_13;
    io_input_13_delay_2 <= io_input_13_delay_1;
    io_input_14_delay_1 <= io_input_14;
  end


endmodule

module TypeB_SkewBuffer (
  input  wire [7:0]    io_input_0,
  input  wire [7:0]    io_input_1,
  input  wire [7:0]    io_input_2,
  input  wire [7:0]    io_input_3,
  input  wire [7:0]    io_input_4,
  input  wire [7:0]    io_input_5,
  input  wire [7:0]    io_input_6,
  input  wire [7:0]    io_input_7,
  input  wire [7:0]    io_input_8,
  input  wire [7:0]    io_input_9,
  input  wire [7:0]    io_input_10,
  input  wire [7:0]    io_input_11,
  input  wire [7:0]    io_input_12,
  input  wire [7:0]    io_input_13,
  input  wire [7:0]    io_input_14,
  input  wire [7:0]    io_input_15,
  output wire [7:0]    io_output_0,
  output wire [7:0]    io_output_1,
  output wire [7:0]    io_output_2,
  output wire [7:0]    io_output_3,
  output wire [7:0]    io_output_4,
  output wire [7:0]    io_output_5,
  output wire [7:0]    io_output_6,
  output wire [7:0]    io_output_7,
  output wire [7:0]    io_output_8,
  output wire [7:0]    io_output_9,
  output wire [7:0]    io_output_10,
  output wire [7:0]    io_output_11,
  output wire [7:0]    io_output_12,
  output wire [7:0]    io_output_13,
  output wire [7:0]    io_output_14,
  output wire [7:0]    io_output_15,
  input  wire          clk,
  input  wire          reset
);

  reg        [7:0]    io_input_0_delay_1;
  reg        [7:0]    io_input_1_delay_1;
  reg        [7:0]    io_input_1_delay_2;
  reg        [7:0]    io_input_2_delay_1;
  reg        [7:0]    io_input_2_delay_2;
  reg        [7:0]    io_input_2_delay_3;
  reg        [7:0]    io_input_3_delay_1;
  reg        [7:0]    io_input_3_delay_2;
  reg        [7:0]    io_input_3_delay_3;
  reg        [7:0]    io_input_3_delay_4;
  reg        [7:0]    io_input_4_delay_1;
  reg        [7:0]    io_input_4_delay_2;
  reg        [7:0]    io_input_4_delay_3;
  reg        [7:0]    io_input_4_delay_4;
  reg        [7:0]    io_input_4_delay_5;
  reg        [7:0]    io_input_5_delay_1;
  reg        [7:0]    io_input_5_delay_2;
  reg        [7:0]    io_input_5_delay_3;
  reg        [7:0]    io_input_5_delay_4;
  reg        [7:0]    io_input_5_delay_5;
  reg        [7:0]    io_input_5_delay_6;
  reg        [7:0]    io_input_6_delay_1;
  reg        [7:0]    io_input_6_delay_2;
  reg        [7:0]    io_input_6_delay_3;
  reg        [7:0]    io_input_6_delay_4;
  reg        [7:0]    io_input_6_delay_5;
  reg        [7:0]    io_input_6_delay_6;
  reg        [7:0]    io_input_6_delay_7;
  reg        [7:0]    io_input_7_delay_1;
  reg        [7:0]    io_input_7_delay_2;
  reg        [7:0]    io_input_7_delay_3;
  reg        [7:0]    io_input_7_delay_4;
  reg        [7:0]    io_input_7_delay_5;
  reg        [7:0]    io_input_7_delay_6;
  reg        [7:0]    io_input_7_delay_7;
  reg        [7:0]    io_input_7_delay_8;
  reg        [7:0]    io_input_8_delay_1;
  reg        [7:0]    io_input_8_delay_2;
  reg        [7:0]    io_input_8_delay_3;
  reg        [7:0]    io_input_8_delay_4;
  reg        [7:0]    io_input_8_delay_5;
  reg        [7:0]    io_input_8_delay_6;
  reg        [7:0]    io_input_8_delay_7;
  reg        [7:0]    io_input_8_delay_8;
  reg        [7:0]    io_input_8_delay_9;
  reg        [7:0]    io_input_9_delay_1;
  reg        [7:0]    io_input_9_delay_2;
  reg        [7:0]    io_input_9_delay_3;
  reg        [7:0]    io_input_9_delay_4;
  reg        [7:0]    io_input_9_delay_5;
  reg        [7:0]    io_input_9_delay_6;
  reg        [7:0]    io_input_9_delay_7;
  reg        [7:0]    io_input_9_delay_8;
  reg        [7:0]    io_input_9_delay_9;
  reg        [7:0]    io_input_9_delay_10;
  reg        [7:0]    io_input_10_delay_1;
  reg        [7:0]    io_input_10_delay_2;
  reg        [7:0]    io_input_10_delay_3;
  reg        [7:0]    io_input_10_delay_4;
  reg        [7:0]    io_input_10_delay_5;
  reg        [7:0]    io_input_10_delay_6;
  reg        [7:0]    io_input_10_delay_7;
  reg        [7:0]    io_input_10_delay_8;
  reg        [7:0]    io_input_10_delay_9;
  reg        [7:0]    io_input_10_delay_10;
  reg        [7:0]    io_input_10_delay_11;
  reg        [7:0]    io_input_11_delay_1;
  reg        [7:0]    io_input_11_delay_2;
  reg        [7:0]    io_input_11_delay_3;
  reg        [7:0]    io_input_11_delay_4;
  reg        [7:0]    io_input_11_delay_5;
  reg        [7:0]    io_input_11_delay_6;
  reg        [7:0]    io_input_11_delay_7;
  reg        [7:0]    io_input_11_delay_8;
  reg        [7:0]    io_input_11_delay_9;
  reg        [7:0]    io_input_11_delay_10;
  reg        [7:0]    io_input_11_delay_11;
  reg        [7:0]    io_input_11_delay_12;
  reg        [7:0]    io_input_12_delay_1;
  reg        [7:0]    io_input_12_delay_2;
  reg        [7:0]    io_input_12_delay_3;
  reg        [7:0]    io_input_12_delay_4;
  reg        [7:0]    io_input_12_delay_5;
  reg        [7:0]    io_input_12_delay_6;
  reg        [7:0]    io_input_12_delay_7;
  reg        [7:0]    io_input_12_delay_8;
  reg        [7:0]    io_input_12_delay_9;
  reg        [7:0]    io_input_12_delay_10;
  reg        [7:0]    io_input_12_delay_11;
  reg        [7:0]    io_input_12_delay_12;
  reg        [7:0]    io_input_12_delay_13;
  reg        [7:0]    io_input_13_delay_1;
  reg        [7:0]    io_input_13_delay_2;
  reg        [7:0]    io_input_13_delay_3;
  reg        [7:0]    io_input_13_delay_4;
  reg        [7:0]    io_input_13_delay_5;
  reg        [7:0]    io_input_13_delay_6;
  reg        [7:0]    io_input_13_delay_7;
  reg        [7:0]    io_input_13_delay_8;
  reg        [7:0]    io_input_13_delay_9;
  reg        [7:0]    io_input_13_delay_10;
  reg        [7:0]    io_input_13_delay_11;
  reg        [7:0]    io_input_13_delay_12;
  reg        [7:0]    io_input_13_delay_13;
  reg        [7:0]    io_input_13_delay_14;
  reg        [7:0]    io_input_14_delay_1;
  reg        [7:0]    io_input_14_delay_2;
  reg        [7:0]    io_input_14_delay_3;
  reg        [7:0]    io_input_14_delay_4;
  reg        [7:0]    io_input_14_delay_5;
  reg        [7:0]    io_input_14_delay_6;
  reg        [7:0]    io_input_14_delay_7;
  reg        [7:0]    io_input_14_delay_8;
  reg        [7:0]    io_input_14_delay_9;
  reg        [7:0]    io_input_14_delay_10;
  reg        [7:0]    io_input_14_delay_11;
  reg        [7:0]    io_input_14_delay_12;
  reg        [7:0]    io_input_14_delay_13;
  reg        [7:0]    io_input_14_delay_14;
  reg        [7:0]    io_input_14_delay_15;
  reg        [7:0]    io_input_15_delay_1;
  reg        [7:0]    io_input_15_delay_2;
  reg        [7:0]    io_input_15_delay_3;
  reg        [7:0]    io_input_15_delay_4;
  reg        [7:0]    io_input_15_delay_5;
  reg        [7:0]    io_input_15_delay_6;
  reg        [7:0]    io_input_15_delay_7;
  reg        [7:0]    io_input_15_delay_8;
  reg        [7:0]    io_input_15_delay_9;
  reg        [7:0]    io_input_15_delay_10;
  reg        [7:0]    io_input_15_delay_11;
  reg        [7:0]    io_input_15_delay_12;
  reg        [7:0]    io_input_15_delay_13;
  reg        [7:0]    io_input_15_delay_14;
  reg        [7:0]    io_input_15_delay_15;
  reg        [7:0]    io_input_15_delay_16;

  assign io_output_0 = io_input_0_delay_1;
  assign io_output_1 = io_input_1_delay_2;
  assign io_output_2 = io_input_2_delay_3;
  assign io_output_3 = io_input_3_delay_4;
  assign io_output_4 = io_input_4_delay_5;
  assign io_output_5 = io_input_5_delay_6;
  assign io_output_6 = io_input_6_delay_7;
  assign io_output_7 = io_input_7_delay_8;
  assign io_output_8 = io_input_8_delay_9;
  assign io_output_9 = io_input_9_delay_10;
  assign io_output_10 = io_input_10_delay_11;
  assign io_output_11 = io_input_11_delay_12;
  assign io_output_12 = io_input_12_delay_13;
  assign io_output_13 = io_input_13_delay_14;
  assign io_output_14 = io_input_14_delay_15;
  assign io_output_15 = io_input_15_delay_16;
  always @(posedge clk) begin
    io_input_0_delay_1 <= io_input_0;
    io_input_1_delay_1 <= io_input_1;
    io_input_1_delay_2 <= io_input_1_delay_1;
    io_input_2_delay_1 <= io_input_2;
    io_input_2_delay_2 <= io_input_2_delay_1;
    io_input_2_delay_3 <= io_input_2_delay_2;
    io_input_3_delay_1 <= io_input_3;
    io_input_3_delay_2 <= io_input_3_delay_1;
    io_input_3_delay_3 <= io_input_3_delay_2;
    io_input_3_delay_4 <= io_input_3_delay_3;
    io_input_4_delay_1 <= io_input_4;
    io_input_4_delay_2 <= io_input_4_delay_1;
    io_input_4_delay_3 <= io_input_4_delay_2;
    io_input_4_delay_4 <= io_input_4_delay_3;
    io_input_4_delay_5 <= io_input_4_delay_4;
    io_input_5_delay_1 <= io_input_5;
    io_input_5_delay_2 <= io_input_5_delay_1;
    io_input_5_delay_3 <= io_input_5_delay_2;
    io_input_5_delay_4 <= io_input_5_delay_3;
    io_input_5_delay_5 <= io_input_5_delay_4;
    io_input_5_delay_6 <= io_input_5_delay_5;
    io_input_6_delay_1 <= io_input_6;
    io_input_6_delay_2 <= io_input_6_delay_1;
    io_input_6_delay_3 <= io_input_6_delay_2;
    io_input_6_delay_4 <= io_input_6_delay_3;
    io_input_6_delay_5 <= io_input_6_delay_4;
    io_input_6_delay_6 <= io_input_6_delay_5;
    io_input_6_delay_7 <= io_input_6_delay_6;
    io_input_7_delay_1 <= io_input_7;
    io_input_7_delay_2 <= io_input_7_delay_1;
    io_input_7_delay_3 <= io_input_7_delay_2;
    io_input_7_delay_4 <= io_input_7_delay_3;
    io_input_7_delay_5 <= io_input_7_delay_4;
    io_input_7_delay_6 <= io_input_7_delay_5;
    io_input_7_delay_7 <= io_input_7_delay_6;
    io_input_7_delay_8 <= io_input_7_delay_7;
    io_input_8_delay_1 <= io_input_8;
    io_input_8_delay_2 <= io_input_8_delay_1;
    io_input_8_delay_3 <= io_input_8_delay_2;
    io_input_8_delay_4 <= io_input_8_delay_3;
    io_input_8_delay_5 <= io_input_8_delay_4;
    io_input_8_delay_6 <= io_input_8_delay_5;
    io_input_8_delay_7 <= io_input_8_delay_6;
    io_input_8_delay_8 <= io_input_8_delay_7;
    io_input_8_delay_9 <= io_input_8_delay_8;
    io_input_9_delay_1 <= io_input_9;
    io_input_9_delay_2 <= io_input_9_delay_1;
    io_input_9_delay_3 <= io_input_9_delay_2;
    io_input_9_delay_4 <= io_input_9_delay_3;
    io_input_9_delay_5 <= io_input_9_delay_4;
    io_input_9_delay_6 <= io_input_9_delay_5;
    io_input_9_delay_7 <= io_input_9_delay_6;
    io_input_9_delay_8 <= io_input_9_delay_7;
    io_input_9_delay_9 <= io_input_9_delay_8;
    io_input_9_delay_10 <= io_input_9_delay_9;
    io_input_10_delay_1 <= io_input_10;
    io_input_10_delay_2 <= io_input_10_delay_1;
    io_input_10_delay_3 <= io_input_10_delay_2;
    io_input_10_delay_4 <= io_input_10_delay_3;
    io_input_10_delay_5 <= io_input_10_delay_4;
    io_input_10_delay_6 <= io_input_10_delay_5;
    io_input_10_delay_7 <= io_input_10_delay_6;
    io_input_10_delay_8 <= io_input_10_delay_7;
    io_input_10_delay_9 <= io_input_10_delay_8;
    io_input_10_delay_10 <= io_input_10_delay_9;
    io_input_10_delay_11 <= io_input_10_delay_10;
    io_input_11_delay_1 <= io_input_11;
    io_input_11_delay_2 <= io_input_11_delay_1;
    io_input_11_delay_3 <= io_input_11_delay_2;
    io_input_11_delay_4 <= io_input_11_delay_3;
    io_input_11_delay_5 <= io_input_11_delay_4;
    io_input_11_delay_6 <= io_input_11_delay_5;
    io_input_11_delay_7 <= io_input_11_delay_6;
    io_input_11_delay_8 <= io_input_11_delay_7;
    io_input_11_delay_9 <= io_input_11_delay_8;
    io_input_11_delay_10 <= io_input_11_delay_9;
    io_input_11_delay_11 <= io_input_11_delay_10;
    io_input_11_delay_12 <= io_input_11_delay_11;
    io_input_12_delay_1 <= io_input_12;
    io_input_12_delay_2 <= io_input_12_delay_1;
    io_input_12_delay_3 <= io_input_12_delay_2;
    io_input_12_delay_4 <= io_input_12_delay_3;
    io_input_12_delay_5 <= io_input_12_delay_4;
    io_input_12_delay_6 <= io_input_12_delay_5;
    io_input_12_delay_7 <= io_input_12_delay_6;
    io_input_12_delay_8 <= io_input_12_delay_7;
    io_input_12_delay_9 <= io_input_12_delay_8;
    io_input_12_delay_10 <= io_input_12_delay_9;
    io_input_12_delay_11 <= io_input_12_delay_10;
    io_input_12_delay_12 <= io_input_12_delay_11;
    io_input_12_delay_13 <= io_input_12_delay_12;
    io_input_13_delay_1 <= io_input_13;
    io_input_13_delay_2 <= io_input_13_delay_1;
    io_input_13_delay_3 <= io_input_13_delay_2;
    io_input_13_delay_4 <= io_input_13_delay_3;
    io_input_13_delay_5 <= io_input_13_delay_4;
    io_input_13_delay_6 <= io_input_13_delay_5;
    io_input_13_delay_7 <= io_input_13_delay_6;
    io_input_13_delay_8 <= io_input_13_delay_7;
    io_input_13_delay_9 <= io_input_13_delay_8;
    io_input_13_delay_10 <= io_input_13_delay_9;
    io_input_13_delay_11 <= io_input_13_delay_10;
    io_input_13_delay_12 <= io_input_13_delay_11;
    io_input_13_delay_13 <= io_input_13_delay_12;
    io_input_13_delay_14 <= io_input_13_delay_13;
    io_input_14_delay_1 <= io_input_14;
    io_input_14_delay_2 <= io_input_14_delay_1;
    io_input_14_delay_3 <= io_input_14_delay_2;
    io_input_14_delay_4 <= io_input_14_delay_3;
    io_input_14_delay_5 <= io_input_14_delay_4;
    io_input_14_delay_6 <= io_input_14_delay_5;
    io_input_14_delay_7 <= io_input_14_delay_6;
    io_input_14_delay_8 <= io_input_14_delay_7;
    io_input_14_delay_9 <= io_input_14_delay_8;
    io_input_14_delay_10 <= io_input_14_delay_9;
    io_input_14_delay_11 <= io_input_14_delay_10;
    io_input_14_delay_12 <= io_input_14_delay_11;
    io_input_14_delay_13 <= io_input_14_delay_12;
    io_input_14_delay_14 <= io_input_14_delay_13;
    io_input_14_delay_15 <= io_input_14_delay_14;
    io_input_15_delay_1 <= io_input_15;
    io_input_15_delay_2 <= io_input_15_delay_1;
    io_input_15_delay_3 <= io_input_15_delay_2;
    io_input_15_delay_4 <= io_input_15_delay_3;
    io_input_15_delay_5 <= io_input_15_delay_4;
    io_input_15_delay_6 <= io_input_15_delay_5;
    io_input_15_delay_7 <= io_input_15_delay_6;
    io_input_15_delay_8 <= io_input_15_delay_7;
    io_input_15_delay_9 <= io_input_15_delay_8;
    io_input_15_delay_10 <= io_input_15_delay_9;
    io_input_15_delay_11 <= io_input_15_delay_10;
    io_input_15_delay_12 <= io_input_15_delay_11;
    io_input_15_delay_13 <= io_input_15_delay_12;
    io_input_15_delay_14 <= io_input_15_delay_13;
    io_input_15_delay_15 <= io_input_15_delay_14;
    io_input_15_delay_16 <= io_input_15_delay_15;
  end


endmodule

module TypeA_SkewBuffer (
  input  wire [7:0]    io_input_0,
  input  wire [7:0]    io_input_1,
  input  wire [7:0]    io_input_2,
  input  wire [7:0]    io_input_3,
  input  wire [7:0]    io_input_4,
  input  wire [7:0]    io_input_5,
  input  wire [7:0]    io_input_6,
  input  wire [7:0]    io_input_7,
  input  wire [7:0]    io_input_8,
  input  wire [7:0]    io_input_9,
  input  wire [7:0]    io_input_10,
  input  wire [7:0]    io_input_11,
  input  wire [7:0]    io_input_12,
  input  wire [7:0]    io_input_13,
  input  wire [7:0]    io_input_14,
  input  wire [7:0]    io_input_15,
  output wire [7:0]    io_output_0,
  output wire [7:0]    io_output_1,
  output wire [7:0]    io_output_2,
  output wire [7:0]    io_output_3,
  output wire [7:0]    io_output_4,
  output wire [7:0]    io_output_5,
  output wire [7:0]    io_output_6,
  output wire [7:0]    io_output_7,
  output wire [7:0]    io_output_8,
  output wire [7:0]    io_output_9,
  output wire [7:0]    io_output_10,
  output wire [7:0]    io_output_11,
  output wire [7:0]    io_output_12,
  output wire [7:0]    io_output_13,
  output wire [7:0]    io_output_14,
  output wire [7:0]    io_output_15,
  input  wire          clk,
  input  wire          reset
);

  reg        [7:0]    io_input_0_delay_1;
  reg        [7:0]    io_input_1_delay_1;
  reg        [7:0]    io_input_1_delay_2;
  reg        [7:0]    io_input_2_delay_1;
  reg        [7:0]    io_input_2_delay_2;
  reg        [7:0]    io_input_2_delay_3;
  reg        [7:0]    io_input_3_delay_1;
  reg        [7:0]    io_input_3_delay_2;
  reg        [7:0]    io_input_3_delay_3;
  reg        [7:0]    io_input_3_delay_4;
  reg        [7:0]    io_input_4_delay_1;
  reg        [7:0]    io_input_4_delay_2;
  reg        [7:0]    io_input_4_delay_3;
  reg        [7:0]    io_input_4_delay_4;
  reg        [7:0]    io_input_4_delay_5;
  reg        [7:0]    io_input_5_delay_1;
  reg        [7:0]    io_input_5_delay_2;
  reg        [7:0]    io_input_5_delay_3;
  reg        [7:0]    io_input_5_delay_4;
  reg        [7:0]    io_input_5_delay_5;
  reg        [7:0]    io_input_5_delay_6;
  reg        [7:0]    io_input_6_delay_1;
  reg        [7:0]    io_input_6_delay_2;
  reg        [7:0]    io_input_6_delay_3;
  reg        [7:0]    io_input_6_delay_4;
  reg        [7:0]    io_input_6_delay_5;
  reg        [7:0]    io_input_6_delay_6;
  reg        [7:0]    io_input_6_delay_7;
  reg        [7:0]    io_input_7_delay_1;
  reg        [7:0]    io_input_7_delay_2;
  reg        [7:0]    io_input_7_delay_3;
  reg        [7:0]    io_input_7_delay_4;
  reg        [7:0]    io_input_7_delay_5;
  reg        [7:0]    io_input_7_delay_6;
  reg        [7:0]    io_input_7_delay_7;
  reg        [7:0]    io_input_7_delay_8;
  reg        [7:0]    io_input_8_delay_1;
  reg        [7:0]    io_input_8_delay_2;
  reg        [7:0]    io_input_8_delay_3;
  reg        [7:0]    io_input_8_delay_4;
  reg        [7:0]    io_input_8_delay_5;
  reg        [7:0]    io_input_8_delay_6;
  reg        [7:0]    io_input_8_delay_7;
  reg        [7:0]    io_input_8_delay_8;
  reg        [7:0]    io_input_8_delay_9;
  reg        [7:0]    io_input_9_delay_1;
  reg        [7:0]    io_input_9_delay_2;
  reg        [7:0]    io_input_9_delay_3;
  reg        [7:0]    io_input_9_delay_4;
  reg        [7:0]    io_input_9_delay_5;
  reg        [7:0]    io_input_9_delay_6;
  reg        [7:0]    io_input_9_delay_7;
  reg        [7:0]    io_input_9_delay_8;
  reg        [7:0]    io_input_9_delay_9;
  reg        [7:0]    io_input_9_delay_10;
  reg        [7:0]    io_input_10_delay_1;
  reg        [7:0]    io_input_10_delay_2;
  reg        [7:0]    io_input_10_delay_3;
  reg        [7:0]    io_input_10_delay_4;
  reg        [7:0]    io_input_10_delay_5;
  reg        [7:0]    io_input_10_delay_6;
  reg        [7:0]    io_input_10_delay_7;
  reg        [7:0]    io_input_10_delay_8;
  reg        [7:0]    io_input_10_delay_9;
  reg        [7:0]    io_input_10_delay_10;
  reg        [7:0]    io_input_10_delay_11;
  reg        [7:0]    io_input_11_delay_1;
  reg        [7:0]    io_input_11_delay_2;
  reg        [7:0]    io_input_11_delay_3;
  reg        [7:0]    io_input_11_delay_4;
  reg        [7:0]    io_input_11_delay_5;
  reg        [7:0]    io_input_11_delay_6;
  reg        [7:0]    io_input_11_delay_7;
  reg        [7:0]    io_input_11_delay_8;
  reg        [7:0]    io_input_11_delay_9;
  reg        [7:0]    io_input_11_delay_10;
  reg        [7:0]    io_input_11_delay_11;
  reg        [7:0]    io_input_11_delay_12;
  reg        [7:0]    io_input_12_delay_1;
  reg        [7:0]    io_input_12_delay_2;
  reg        [7:0]    io_input_12_delay_3;
  reg        [7:0]    io_input_12_delay_4;
  reg        [7:0]    io_input_12_delay_5;
  reg        [7:0]    io_input_12_delay_6;
  reg        [7:0]    io_input_12_delay_7;
  reg        [7:0]    io_input_12_delay_8;
  reg        [7:0]    io_input_12_delay_9;
  reg        [7:0]    io_input_12_delay_10;
  reg        [7:0]    io_input_12_delay_11;
  reg        [7:0]    io_input_12_delay_12;
  reg        [7:0]    io_input_12_delay_13;
  reg        [7:0]    io_input_13_delay_1;
  reg        [7:0]    io_input_13_delay_2;
  reg        [7:0]    io_input_13_delay_3;
  reg        [7:0]    io_input_13_delay_4;
  reg        [7:0]    io_input_13_delay_5;
  reg        [7:0]    io_input_13_delay_6;
  reg        [7:0]    io_input_13_delay_7;
  reg        [7:0]    io_input_13_delay_8;
  reg        [7:0]    io_input_13_delay_9;
  reg        [7:0]    io_input_13_delay_10;
  reg        [7:0]    io_input_13_delay_11;
  reg        [7:0]    io_input_13_delay_12;
  reg        [7:0]    io_input_13_delay_13;
  reg        [7:0]    io_input_13_delay_14;
  reg        [7:0]    io_input_14_delay_1;
  reg        [7:0]    io_input_14_delay_2;
  reg        [7:0]    io_input_14_delay_3;
  reg        [7:0]    io_input_14_delay_4;
  reg        [7:0]    io_input_14_delay_5;
  reg        [7:0]    io_input_14_delay_6;
  reg        [7:0]    io_input_14_delay_7;
  reg        [7:0]    io_input_14_delay_8;
  reg        [7:0]    io_input_14_delay_9;
  reg        [7:0]    io_input_14_delay_10;
  reg        [7:0]    io_input_14_delay_11;
  reg        [7:0]    io_input_14_delay_12;
  reg        [7:0]    io_input_14_delay_13;
  reg        [7:0]    io_input_14_delay_14;
  reg        [7:0]    io_input_14_delay_15;
  reg        [7:0]    io_input_15_delay_1;
  reg        [7:0]    io_input_15_delay_2;
  reg        [7:0]    io_input_15_delay_3;
  reg        [7:0]    io_input_15_delay_4;
  reg        [7:0]    io_input_15_delay_5;
  reg        [7:0]    io_input_15_delay_6;
  reg        [7:0]    io_input_15_delay_7;
  reg        [7:0]    io_input_15_delay_8;
  reg        [7:0]    io_input_15_delay_9;
  reg        [7:0]    io_input_15_delay_10;
  reg        [7:0]    io_input_15_delay_11;
  reg        [7:0]    io_input_15_delay_12;
  reg        [7:0]    io_input_15_delay_13;
  reg        [7:0]    io_input_15_delay_14;
  reg        [7:0]    io_input_15_delay_15;
  reg        [7:0]    io_input_15_delay_16;

  assign io_output_0 = io_input_0_delay_1;
  assign io_output_1 = io_input_1_delay_2;
  assign io_output_2 = io_input_2_delay_3;
  assign io_output_3 = io_input_3_delay_4;
  assign io_output_4 = io_input_4_delay_5;
  assign io_output_5 = io_input_5_delay_6;
  assign io_output_6 = io_input_6_delay_7;
  assign io_output_7 = io_input_7_delay_8;
  assign io_output_8 = io_input_8_delay_9;
  assign io_output_9 = io_input_9_delay_10;
  assign io_output_10 = io_input_10_delay_11;
  assign io_output_11 = io_input_11_delay_12;
  assign io_output_12 = io_input_12_delay_13;
  assign io_output_13 = io_input_13_delay_14;
  assign io_output_14 = io_input_14_delay_15;
  assign io_output_15 = io_input_15_delay_16;
  always @(posedge clk) begin
    io_input_0_delay_1 <= io_input_0;
    io_input_1_delay_1 <= io_input_1;
    io_input_1_delay_2 <= io_input_1_delay_1;
    io_input_2_delay_1 <= io_input_2;
    io_input_2_delay_2 <= io_input_2_delay_1;
    io_input_2_delay_3 <= io_input_2_delay_2;
    io_input_3_delay_1 <= io_input_3;
    io_input_3_delay_2 <= io_input_3_delay_1;
    io_input_3_delay_3 <= io_input_3_delay_2;
    io_input_3_delay_4 <= io_input_3_delay_3;
    io_input_4_delay_1 <= io_input_4;
    io_input_4_delay_2 <= io_input_4_delay_1;
    io_input_4_delay_3 <= io_input_4_delay_2;
    io_input_4_delay_4 <= io_input_4_delay_3;
    io_input_4_delay_5 <= io_input_4_delay_4;
    io_input_5_delay_1 <= io_input_5;
    io_input_5_delay_2 <= io_input_5_delay_1;
    io_input_5_delay_3 <= io_input_5_delay_2;
    io_input_5_delay_4 <= io_input_5_delay_3;
    io_input_5_delay_5 <= io_input_5_delay_4;
    io_input_5_delay_6 <= io_input_5_delay_5;
    io_input_6_delay_1 <= io_input_6;
    io_input_6_delay_2 <= io_input_6_delay_1;
    io_input_6_delay_3 <= io_input_6_delay_2;
    io_input_6_delay_4 <= io_input_6_delay_3;
    io_input_6_delay_5 <= io_input_6_delay_4;
    io_input_6_delay_6 <= io_input_6_delay_5;
    io_input_6_delay_7 <= io_input_6_delay_6;
    io_input_7_delay_1 <= io_input_7;
    io_input_7_delay_2 <= io_input_7_delay_1;
    io_input_7_delay_3 <= io_input_7_delay_2;
    io_input_7_delay_4 <= io_input_7_delay_3;
    io_input_7_delay_5 <= io_input_7_delay_4;
    io_input_7_delay_6 <= io_input_7_delay_5;
    io_input_7_delay_7 <= io_input_7_delay_6;
    io_input_7_delay_8 <= io_input_7_delay_7;
    io_input_8_delay_1 <= io_input_8;
    io_input_8_delay_2 <= io_input_8_delay_1;
    io_input_8_delay_3 <= io_input_8_delay_2;
    io_input_8_delay_4 <= io_input_8_delay_3;
    io_input_8_delay_5 <= io_input_8_delay_4;
    io_input_8_delay_6 <= io_input_8_delay_5;
    io_input_8_delay_7 <= io_input_8_delay_6;
    io_input_8_delay_8 <= io_input_8_delay_7;
    io_input_8_delay_9 <= io_input_8_delay_8;
    io_input_9_delay_1 <= io_input_9;
    io_input_9_delay_2 <= io_input_9_delay_1;
    io_input_9_delay_3 <= io_input_9_delay_2;
    io_input_9_delay_4 <= io_input_9_delay_3;
    io_input_9_delay_5 <= io_input_9_delay_4;
    io_input_9_delay_6 <= io_input_9_delay_5;
    io_input_9_delay_7 <= io_input_9_delay_6;
    io_input_9_delay_8 <= io_input_9_delay_7;
    io_input_9_delay_9 <= io_input_9_delay_8;
    io_input_9_delay_10 <= io_input_9_delay_9;
    io_input_10_delay_1 <= io_input_10;
    io_input_10_delay_2 <= io_input_10_delay_1;
    io_input_10_delay_3 <= io_input_10_delay_2;
    io_input_10_delay_4 <= io_input_10_delay_3;
    io_input_10_delay_5 <= io_input_10_delay_4;
    io_input_10_delay_6 <= io_input_10_delay_5;
    io_input_10_delay_7 <= io_input_10_delay_6;
    io_input_10_delay_8 <= io_input_10_delay_7;
    io_input_10_delay_9 <= io_input_10_delay_8;
    io_input_10_delay_10 <= io_input_10_delay_9;
    io_input_10_delay_11 <= io_input_10_delay_10;
    io_input_11_delay_1 <= io_input_11;
    io_input_11_delay_2 <= io_input_11_delay_1;
    io_input_11_delay_3 <= io_input_11_delay_2;
    io_input_11_delay_4 <= io_input_11_delay_3;
    io_input_11_delay_5 <= io_input_11_delay_4;
    io_input_11_delay_6 <= io_input_11_delay_5;
    io_input_11_delay_7 <= io_input_11_delay_6;
    io_input_11_delay_8 <= io_input_11_delay_7;
    io_input_11_delay_9 <= io_input_11_delay_8;
    io_input_11_delay_10 <= io_input_11_delay_9;
    io_input_11_delay_11 <= io_input_11_delay_10;
    io_input_11_delay_12 <= io_input_11_delay_11;
    io_input_12_delay_1 <= io_input_12;
    io_input_12_delay_2 <= io_input_12_delay_1;
    io_input_12_delay_3 <= io_input_12_delay_2;
    io_input_12_delay_4 <= io_input_12_delay_3;
    io_input_12_delay_5 <= io_input_12_delay_4;
    io_input_12_delay_6 <= io_input_12_delay_5;
    io_input_12_delay_7 <= io_input_12_delay_6;
    io_input_12_delay_8 <= io_input_12_delay_7;
    io_input_12_delay_9 <= io_input_12_delay_8;
    io_input_12_delay_10 <= io_input_12_delay_9;
    io_input_12_delay_11 <= io_input_12_delay_10;
    io_input_12_delay_12 <= io_input_12_delay_11;
    io_input_12_delay_13 <= io_input_12_delay_12;
    io_input_13_delay_1 <= io_input_13;
    io_input_13_delay_2 <= io_input_13_delay_1;
    io_input_13_delay_3 <= io_input_13_delay_2;
    io_input_13_delay_4 <= io_input_13_delay_3;
    io_input_13_delay_5 <= io_input_13_delay_4;
    io_input_13_delay_6 <= io_input_13_delay_5;
    io_input_13_delay_7 <= io_input_13_delay_6;
    io_input_13_delay_8 <= io_input_13_delay_7;
    io_input_13_delay_9 <= io_input_13_delay_8;
    io_input_13_delay_10 <= io_input_13_delay_9;
    io_input_13_delay_11 <= io_input_13_delay_10;
    io_input_13_delay_12 <= io_input_13_delay_11;
    io_input_13_delay_13 <= io_input_13_delay_12;
    io_input_13_delay_14 <= io_input_13_delay_13;
    io_input_14_delay_1 <= io_input_14;
    io_input_14_delay_2 <= io_input_14_delay_1;
    io_input_14_delay_3 <= io_input_14_delay_2;
    io_input_14_delay_4 <= io_input_14_delay_3;
    io_input_14_delay_5 <= io_input_14_delay_4;
    io_input_14_delay_6 <= io_input_14_delay_5;
    io_input_14_delay_7 <= io_input_14_delay_6;
    io_input_14_delay_8 <= io_input_14_delay_7;
    io_input_14_delay_9 <= io_input_14_delay_8;
    io_input_14_delay_10 <= io_input_14_delay_9;
    io_input_14_delay_11 <= io_input_14_delay_10;
    io_input_14_delay_12 <= io_input_14_delay_11;
    io_input_14_delay_13 <= io_input_14_delay_12;
    io_input_14_delay_14 <= io_input_14_delay_13;
    io_input_14_delay_15 <= io_input_14_delay_14;
    io_input_15_delay_1 <= io_input_15;
    io_input_15_delay_2 <= io_input_15_delay_1;
    io_input_15_delay_3 <= io_input_15_delay_2;
    io_input_15_delay_4 <= io_input_15_delay_3;
    io_input_15_delay_5 <= io_input_15_delay_4;
    io_input_15_delay_6 <= io_input_15_delay_5;
    io_input_15_delay_7 <= io_input_15_delay_6;
    io_input_15_delay_8 <= io_input_15_delay_7;
    io_input_15_delay_9 <= io_input_15_delay_8;
    io_input_15_delay_10 <= io_input_15_delay_9;
    io_input_15_delay_11 <= io_input_15_delay_10;
    io_input_15_delay_12 <= io_input_15_delay_11;
    io_input_15_delay_13 <= io_input_15_delay_12;
    io_input_15_delay_14 <= io_input_15_delay_13;
    io_input_15_delay_15 <= io_input_15_delay_14;
    io_input_15_delay_16 <= io_input_15_delay_15;
  end


endmodule

module ProcessingElement_255 (
  input  wire [7:0]    io_inputA,
  input  wire [7:0]    io_inputB,
  input  wire          io_outputCaptureEnableC,
  input  wire          io_resetPartialC,
  output wire [25:0]   io_outputC,
  input  wire          clk,
  input  wire          reset
);

  wire       [25:0]   _zz__zz_io_outputC_1;
  wire       [25:0]   _zz__zz_io_outputC_1_1;
  wire       [25:0]   _zz__zz_io_outputC_1_2;
  wire       [15:0]   _zz_io_outputC;
  reg        [25:0]   _zz_io_outputC_1;

  assign _zz__zz_io_outputC_1 = {{10{_zz_io_outputC[15]}}, _zz_io_outputC};
  assign _zz__zz_io_outputC_1_1 = ($signed(_zz__zz_io_outputC_1_2) + $signed(_zz_io_outputC_1));
  assign _zz__zz_io_outputC_1_2 = {{10{_zz_io_outputC[15]}}, _zz_io_outputC};
  assign _zz_io_outputC = ($signed(io_inputA) * $signed(io_inputB));
  assign io_outputC = _zz_io_outputC_1;
  always @(posedge clk) begin
    if(reset) begin
      _zz_io_outputC_1 <= 26'h0;
    end else begin
      _zz_io_outputC_1 <= (io_resetPartialC ? _zz__zz_io_outputC_1 : _zz__zz_io_outputC_1_1);
    end
  end


endmodule

//ProcessingElement_254 replaced by ProcessingElement_240

//ProcessingElement_253 replaced by ProcessingElement_240

//ProcessingElement_252 replaced by ProcessingElement_240

//ProcessingElement_251 replaced by ProcessingElement_240

//ProcessingElement_250 replaced by ProcessingElement_240

//ProcessingElement_249 replaced by ProcessingElement_240

//ProcessingElement_248 replaced by ProcessingElement_240

//ProcessingElement_247 replaced by ProcessingElement_240

//ProcessingElement_246 replaced by ProcessingElement_240

//ProcessingElement_245 replaced by ProcessingElement_240

//ProcessingElement_244 replaced by ProcessingElement_240

//ProcessingElement_243 replaced by ProcessingElement_240

//ProcessingElement_242 replaced by ProcessingElement_240

//ProcessingElement_241 replaced by ProcessingElement_240

module ProcessingElement_240 (
  input  wire [7:0]    io_inputA,
  input  wire [7:0]    io_inputB,
  input  wire [25:0]   io_inputC,
  input  wire          io_outputCaptureEnableC,
  input  wire          io_resetPartialC,
  output wire [7:0]    io_outputA,
  output wire [25:0]   io_outputC,
  input  wire          clk,
  input  wire          reset
);

  wire       [25:0]   _zz__zz_io_outputC_1;
  wire       [25:0]   _zz__zz_io_outputC_1_1;
  wire       [25:0]   _zz__zz_io_outputC_1_2;
  reg        [7:0]    io_inputA_regNext;
  wire       [15:0]   _zz_io_outputC;
  reg        [25:0]   _zz_io_outputC_1;
  reg        [25:0]   _zz_io_outputC_2;

  assign _zz__zz_io_outputC_1 = {{10{_zz_io_outputC[15]}}, _zz_io_outputC};
  assign _zz__zz_io_outputC_1_1 = ($signed(_zz__zz_io_outputC_1_2) + $signed(_zz_io_outputC_1));
  assign _zz__zz_io_outputC_1_2 = {{10{_zz_io_outputC[15]}}, _zz_io_outputC};
  assign io_outputA = io_inputA_regNext;
  assign _zz_io_outputC = ($signed(io_inputA) * $signed(io_inputB));
  assign io_outputC = _zz_io_outputC_2;
  always @(posedge clk) begin
    if(reset) begin
      io_inputA_regNext <= 8'h0;
      _zz_io_outputC_1 <= 26'h0;
      _zz_io_outputC_2 <= 26'h0;
    end else begin
      io_inputA_regNext <= io_inputA;
      _zz_io_outputC_1 <= (io_resetPartialC ? _zz__zz_io_outputC_1 : _zz__zz_io_outputC_1_1);
      _zz_io_outputC_2 <= (io_outputCaptureEnableC ? _zz_io_outputC_1 : io_inputC);
    end
  end


endmodule

//ProcessingElement_239 replaced by ProcessingElement_15

//ProcessingElement_238 replaced by ProcessingElement_16

//ProcessingElement_237 replaced by ProcessingElement_16

//ProcessingElement_236 replaced by ProcessingElement_16

//ProcessingElement_235 replaced by ProcessingElement_16

//ProcessingElement_234 replaced by ProcessingElement_16

//ProcessingElement_233 replaced by ProcessingElement_16

//ProcessingElement_232 replaced by ProcessingElement_16

//ProcessingElement_231 replaced by ProcessingElement_16

//ProcessingElement_230 replaced by ProcessingElement_16

//ProcessingElement_229 replaced by ProcessingElement_16

//ProcessingElement_228 replaced by ProcessingElement_16

//ProcessingElement_227 replaced by ProcessingElement_16

//ProcessingElement_226 replaced by ProcessingElement_16

//ProcessingElement_225 replaced by ProcessingElement_16

//ProcessingElement_224 replaced by ProcessingElement_16

//ProcessingElement_223 replaced by ProcessingElement_15

//ProcessingElement_222 replaced by ProcessingElement_16

//ProcessingElement_221 replaced by ProcessingElement_16

//ProcessingElement_220 replaced by ProcessingElement_16

//ProcessingElement_219 replaced by ProcessingElement_16

//ProcessingElement_218 replaced by ProcessingElement_16

//ProcessingElement_217 replaced by ProcessingElement_16

//ProcessingElement_216 replaced by ProcessingElement_16

//ProcessingElement_215 replaced by ProcessingElement_16

//ProcessingElement_214 replaced by ProcessingElement_16

//ProcessingElement_213 replaced by ProcessingElement_16

//ProcessingElement_212 replaced by ProcessingElement_16

//ProcessingElement_211 replaced by ProcessingElement_16

//ProcessingElement_210 replaced by ProcessingElement_16

//ProcessingElement_209 replaced by ProcessingElement_16

//ProcessingElement_208 replaced by ProcessingElement_16

//ProcessingElement_207 replaced by ProcessingElement_15

//ProcessingElement_206 replaced by ProcessingElement_16

//ProcessingElement_205 replaced by ProcessingElement_16

//ProcessingElement_204 replaced by ProcessingElement_16

//ProcessingElement_203 replaced by ProcessingElement_16

//ProcessingElement_202 replaced by ProcessingElement_16

//ProcessingElement_201 replaced by ProcessingElement_16

//ProcessingElement_200 replaced by ProcessingElement_16

//ProcessingElement_199 replaced by ProcessingElement_16

//ProcessingElement_198 replaced by ProcessingElement_16

//ProcessingElement_197 replaced by ProcessingElement_16

//ProcessingElement_196 replaced by ProcessingElement_16

//ProcessingElement_195 replaced by ProcessingElement_16

//ProcessingElement_194 replaced by ProcessingElement_16

//ProcessingElement_193 replaced by ProcessingElement_16

//ProcessingElement_192 replaced by ProcessingElement_16

//ProcessingElement_191 replaced by ProcessingElement_15

//ProcessingElement_190 replaced by ProcessingElement_16

//ProcessingElement_189 replaced by ProcessingElement_16

//ProcessingElement_188 replaced by ProcessingElement_16

//ProcessingElement_187 replaced by ProcessingElement_16

//ProcessingElement_186 replaced by ProcessingElement_16

//ProcessingElement_185 replaced by ProcessingElement_16

//ProcessingElement_184 replaced by ProcessingElement_16

//ProcessingElement_183 replaced by ProcessingElement_16

//ProcessingElement_182 replaced by ProcessingElement_16

//ProcessingElement_181 replaced by ProcessingElement_16

//ProcessingElement_180 replaced by ProcessingElement_16

//ProcessingElement_179 replaced by ProcessingElement_16

//ProcessingElement_178 replaced by ProcessingElement_16

//ProcessingElement_177 replaced by ProcessingElement_16

//ProcessingElement_176 replaced by ProcessingElement_16

//ProcessingElement_175 replaced by ProcessingElement_15

//ProcessingElement_174 replaced by ProcessingElement_16

//ProcessingElement_173 replaced by ProcessingElement_16

//ProcessingElement_172 replaced by ProcessingElement_16

//ProcessingElement_171 replaced by ProcessingElement_16

//ProcessingElement_170 replaced by ProcessingElement_16

//ProcessingElement_169 replaced by ProcessingElement_16

//ProcessingElement_168 replaced by ProcessingElement_16

//ProcessingElement_167 replaced by ProcessingElement_16

//ProcessingElement_166 replaced by ProcessingElement_16

//ProcessingElement_165 replaced by ProcessingElement_16

//ProcessingElement_164 replaced by ProcessingElement_16

//ProcessingElement_163 replaced by ProcessingElement_16

//ProcessingElement_162 replaced by ProcessingElement_16

//ProcessingElement_161 replaced by ProcessingElement_16

//ProcessingElement_160 replaced by ProcessingElement_16

//ProcessingElement_159 replaced by ProcessingElement_15

//ProcessingElement_158 replaced by ProcessingElement_16

//ProcessingElement_157 replaced by ProcessingElement_16

//ProcessingElement_156 replaced by ProcessingElement_16

//ProcessingElement_155 replaced by ProcessingElement_16

//ProcessingElement_154 replaced by ProcessingElement_16

//ProcessingElement_153 replaced by ProcessingElement_16

//ProcessingElement_152 replaced by ProcessingElement_16

//ProcessingElement_151 replaced by ProcessingElement_16

//ProcessingElement_150 replaced by ProcessingElement_16

//ProcessingElement_149 replaced by ProcessingElement_16

//ProcessingElement_148 replaced by ProcessingElement_16

//ProcessingElement_147 replaced by ProcessingElement_16

//ProcessingElement_146 replaced by ProcessingElement_16

//ProcessingElement_145 replaced by ProcessingElement_16

//ProcessingElement_144 replaced by ProcessingElement_16

//ProcessingElement_143 replaced by ProcessingElement_15

//ProcessingElement_142 replaced by ProcessingElement_16

//ProcessingElement_141 replaced by ProcessingElement_16

//ProcessingElement_140 replaced by ProcessingElement_16

//ProcessingElement_139 replaced by ProcessingElement_16

//ProcessingElement_138 replaced by ProcessingElement_16

//ProcessingElement_137 replaced by ProcessingElement_16

//ProcessingElement_136 replaced by ProcessingElement_16

//ProcessingElement_135 replaced by ProcessingElement_16

//ProcessingElement_134 replaced by ProcessingElement_16

//ProcessingElement_133 replaced by ProcessingElement_16

//ProcessingElement_132 replaced by ProcessingElement_16

//ProcessingElement_131 replaced by ProcessingElement_16

//ProcessingElement_130 replaced by ProcessingElement_16

//ProcessingElement_129 replaced by ProcessingElement_16

//ProcessingElement_128 replaced by ProcessingElement_16

//ProcessingElement_127 replaced by ProcessingElement_15

//ProcessingElement_126 replaced by ProcessingElement_16

//ProcessingElement_125 replaced by ProcessingElement_16

//ProcessingElement_124 replaced by ProcessingElement_16

//ProcessingElement_123 replaced by ProcessingElement_16

//ProcessingElement_122 replaced by ProcessingElement_16

//ProcessingElement_121 replaced by ProcessingElement_16

//ProcessingElement_120 replaced by ProcessingElement_16

//ProcessingElement_119 replaced by ProcessingElement_16

//ProcessingElement_118 replaced by ProcessingElement_16

//ProcessingElement_117 replaced by ProcessingElement_16

//ProcessingElement_116 replaced by ProcessingElement_16

//ProcessingElement_115 replaced by ProcessingElement_16

//ProcessingElement_114 replaced by ProcessingElement_16

//ProcessingElement_113 replaced by ProcessingElement_16

//ProcessingElement_112 replaced by ProcessingElement_16

//ProcessingElement_111 replaced by ProcessingElement_15

//ProcessingElement_110 replaced by ProcessingElement_16

//ProcessingElement_109 replaced by ProcessingElement_16

//ProcessingElement_108 replaced by ProcessingElement_16

//ProcessingElement_107 replaced by ProcessingElement_16

//ProcessingElement_106 replaced by ProcessingElement_16

//ProcessingElement_105 replaced by ProcessingElement_16

//ProcessingElement_104 replaced by ProcessingElement_16

//ProcessingElement_103 replaced by ProcessingElement_16

//ProcessingElement_102 replaced by ProcessingElement_16

//ProcessingElement_101 replaced by ProcessingElement_16

//ProcessingElement_100 replaced by ProcessingElement_16

//ProcessingElement_99 replaced by ProcessingElement_16

//ProcessingElement_98 replaced by ProcessingElement_16

//ProcessingElement_97 replaced by ProcessingElement_16

//ProcessingElement_96 replaced by ProcessingElement_16

//ProcessingElement_95 replaced by ProcessingElement_15

//ProcessingElement_94 replaced by ProcessingElement_16

//ProcessingElement_93 replaced by ProcessingElement_16

//ProcessingElement_92 replaced by ProcessingElement_16

//ProcessingElement_91 replaced by ProcessingElement_16

//ProcessingElement_90 replaced by ProcessingElement_16

//ProcessingElement_89 replaced by ProcessingElement_16

//ProcessingElement_88 replaced by ProcessingElement_16

//ProcessingElement_87 replaced by ProcessingElement_16

//ProcessingElement_86 replaced by ProcessingElement_16

//ProcessingElement_85 replaced by ProcessingElement_16

//ProcessingElement_84 replaced by ProcessingElement_16

//ProcessingElement_83 replaced by ProcessingElement_16

//ProcessingElement_82 replaced by ProcessingElement_16

//ProcessingElement_81 replaced by ProcessingElement_16

//ProcessingElement_80 replaced by ProcessingElement_16

//ProcessingElement_79 replaced by ProcessingElement_15

//ProcessingElement_78 replaced by ProcessingElement_16

//ProcessingElement_77 replaced by ProcessingElement_16

//ProcessingElement_76 replaced by ProcessingElement_16

//ProcessingElement_75 replaced by ProcessingElement_16

//ProcessingElement_74 replaced by ProcessingElement_16

//ProcessingElement_73 replaced by ProcessingElement_16

//ProcessingElement_72 replaced by ProcessingElement_16

//ProcessingElement_71 replaced by ProcessingElement_16

//ProcessingElement_70 replaced by ProcessingElement_16

//ProcessingElement_69 replaced by ProcessingElement_16

//ProcessingElement_68 replaced by ProcessingElement_16

//ProcessingElement_67 replaced by ProcessingElement_16

//ProcessingElement_66 replaced by ProcessingElement_16

//ProcessingElement_65 replaced by ProcessingElement_16

//ProcessingElement_64 replaced by ProcessingElement_16

//ProcessingElement_63 replaced by ProcessingElement_15

//ProcessingElement_62 replaced by ProcessingElement_16

//ProcessingElement_61 replaced by ProcessingElement_16

//ProcessingElement_60 replaced by ProcessingElement_16

//ProcessingElement_59 replaced by ProcessingElement_16

//ProcessingElement_58 replaced by ProcessingElement_16

//ProcessingElement_57 replaced by ProcessingElement_16

//ProcessingElement_56 replaced by ProcessingElement_16

//ProcessingElement_55 replaced by ProcessingElement_16

//ProcessingElement_54 replaced by ProcessingElement_16

//ProcessingElement_53 replaced by ProcessingElement_16

//ProcessingElement_52 replaced by ProcessingElement_16

//ProcessingElement_51 replaced by ProcessingElement_16

//ProcessingElement_50 replaced by ProcessingElement_16

//ProcessingElement_49 replaced by ProcessingElement_16

//ProcessingElement_48 replaced by ProcessingElement_16

//ProcessingElement_47 replaced by ProcessingElement_15

//ProcessingElement_46 replaced by ProcessingElement_16

//ProcessingElement_45 replaced by ProcessingElement_16

//ProcessingElement_44 replaced by ProcessingElement_16

//ProcessingElement_43 replaced by ProcessingElement_16

//ProcessingElement_42 replaced by ProcessingElement_16

//ProcessingElement_41 replaced by ProcessingElement_16

//ProcessingElement_40 replaced by ProcessingElement_16

//ProcessingElement_39 replaced by ProcessingElement_16

//ProcessingElement_38 replaced by ProcessingElement_16

//ProcessingElement_37 replaced by ProcessingElement_16

//ProcessingElement_36 replaced by ProcessingElement_16

//ProcessingElement_35 replaced by ProcessingElement_16

//ProcessingElement_34 replaced by ProcessingElement_16

//ProcessingElement_33 replaced by ProcessingElement_16

//ProcessingElement_32 replaced by ProcessingElement_16

//ProcessingElement_31 replaced by ProcessingElement_15

//ProcessingElement_30 replaced by ProcessingElement_16

//ProcessingElement_29 replaced by ProcessingElement_16

//ProcessingElement_28 replaced by ProcessingElement_16

//ProcessingElement_27 replaced by ProcessingElement_16

//ProcessingElement_26 replaced by ProcessingElement_16

//ProcessingElement_25 replaced by ProcessingElement_16

//ProcessingElement_24 replaced by ProcessingElement_16

//ProcessingElement_23 replaced by ProcessingElement_16

//ProcessingElement_22 replaced by ProcessingElement_16

//ProcessingElement_21 replaced by ProcessingElement_16

//ProcessingElement_20 replaced by ProcessingElement_16

//ProcessingElement_19 replaced by ProcessingElement_16

//ProcessingElement_18 replaced by ProcessingElement_16

//ProcessingElement_17 replaced by ProcessingElement_16

module ProcessingElement_16 (
  input  wire [7:0]    io_inputA,
  input  wire [7:0]    io_inputB,
  input  wire [25:0]   io_inputC,
  input  wire          io_outputCaptureEnableC,
  input  wire          io_resetPartialC,
  output wire [7:0]    io_outputA,
  output wire [7:0]    io_outputB,
  output wire [25:0]   io_outputC,
  input  wire          clk,
  input  wire          reset
);

  wire       [25:0]   _zz__zz_io_outputC_1;   // sign extension
  wire       [25:0]   _zz__zz_io_outputC_1_1; // current matmul + past matmul(_zz_io_outputC_1)
  wire       [25:0]   _zz__zz_io_outputC_1_2; // sign extension
  reg        [7:0]    io_inputA_regNext;
  reg        [7:0]    io_inputB_regNext;
  wire       [15:0]   _zz_io_outputC;         // MatMul result
  reg        [25:0]   _zz_io_outputC_1;       // past matmul accumulated
  reg        [25:0]   _zz_io_outputC_2;       // current matmul or bypass io_outputC

  assign _zz__zz_io_outputC_1 = {{10{_zz_io_outputC[15]}}, _zz_io_outputC};
  assign _zz__zz_io_outputC_1_1 = ($signed(_zz__zz_io_outputC_1_2) + $signed(_zz_io_outputC_1));
  assign _zz__zz_io_outputC_1_2 = {{10{_zz_io_outputC[15]}}, _zz_io_outputC};
  assign io_outputA = io_inputA_regNext;
  assign io_outputB = io_inputB_regNext;
  assign _zz_io_outputC = ($signed(io_inputA) * $signed(io_inputB));
  assign io_outputC = _zz_io_outputC_2;
  always @(posedge clk) begin
    if(reset) begin
      io_inputA_regNext <= 8'h0;
      io_inputB_regNext <= 8'h0;
      _zz_io_outputC_1 <= 26'h0;
      _zz_io_outputC_2 <= 26'h0;
    end else begin
      io_inputA_regNext <= io_inputA;
      io_inputB_regNext <= io_inputB;
      _zz_io_outputC_1 <= (io_resetPartialC ? _zz__zz_io_outputC_1 : _zz__zz_io_outputC_1_1);
      _zz_io_outputC_2 <= (io_outputCaptureEnableC ? _zz_io_outputC_1 : io_inputC);
    end
  end


endmodule

module ProcessingElement_15 (
  input  wire [7:0]    io_inputA,
  input  wire [7:0]    io_inputB,
  input  wire          io_outputCaptureEnableC,
  input  wire          io_resetPartialC,
  output wire [7:0]    io_outputB,
  output wire [25:0]   io_outputC,
  input  wire          clk,
  input  wire          reset
);

  wire       [25:0]   _zz__zz_io_outputC_1;
  wire       [25:0]   _zz__zz_io_outputC_1_1;
  wire       [25:0]   _zz__zz_io_outputC_1_2;
  reg        [7:0]    io_inputB_regNext;
  wire       [15:0]   _zz_io_outputC;
  reg        [25:0]   _zz_io_outputC_1;

  assign _zz__zz_io_outputC_1 = {{10{_zz_io_outputC[15]}}, _zz_io_outputC};
  assign _zz__zz_io_outputC_1_1 = ($signed(_zz__zz_io_outputC_1_2) + $signed(_zz_io_outputC_1));
  assign _zz__zz_io_outputC_1_2 = {{10{_zz_io_outputC[15]}}, _zz_io_outputC};
  assign io_outputB = io_inputB_regNext;
  assign _zz_io_outputC = ($signed(io_inputA) * $signed(io_inputB));
  assign io_outputC = _zz_io_outputC_1;
  always @(posedge clk) begin
    if(reset) begin
      io_inputB_regNext <= 8'h0;
      _zz_io_outputC_1 <= 26'h0;
    end else begin
      io_inputB_regNext <= io_inputB;
      _zz_io_outputC_1 <= (io_resetPartialC ? _zz__zz_io_outputC_1 : _zz__zz_io_outputC_1_1);
    end
  end


endmodule

//ProcessingElement_14 replaced by ProcessingElement

//ProcessingElement_13 replaced by ProcessingElement

//ProcessingElement_12 replaced by ProcessingElement

//ProcessingElement_11 replaced by ProcessingElement

//ProcessingElement_10 replaced by ProcessingElement

//ProcessingElement_9 replaced by ProcessingElement

//ProcessingElement_8 replaced by ProcessingElement

//ProcessingElement_7 replaced by ProcessingElement

//ProcessingElement_6 replaced by ProcessingElement

//ProcessingElement_5 replaced by ProcessingElement

//ProcessingElement_4 replaced by ProcessingElement

//ProcessingElement_3 replaced by ProcessingElement

//ProcessingElement_2 replaced by ProcessingElement

//ProcessingElement_1 replaced by ProcessingElement

module ProcessingElement (
  input  wire [7:0]    io_inputA,
  input  wire [7:0]    io_inputB,
  input  wire          io_outputCaptureEnableC,
  input  wire          io_resetPartialC,
  output wire [7:0]    io_outputA,
  output wire [7:0]    io_outputB,
  output wire [25:0]   io_outputC,
  input  wire          clk,
  input  wire          reset
);

  wire       [25:0]   _zz__zz_io_outputC_1;
  wire       [25:0]   _zz__zz_io_outputC_1_1;
  wire       [25:0]   _zz__zz_io_outputC_1_2;
  reg        [7:0]    io_inputA_regNext;
  reg        [7:0]    io_inputB_regNext;
  wire       [15:0]   _zz_io_outputC;
  reg        [25:0]   _zz_io_outputC_1;

  assign _zz__zz_io_outputC_1 = {{10{_zz_io_outputC[15]}}, _zz_io_outputC};
  assign _zz__zz_io_outputC_1_1 = ($signed(_zz__zz_io_outputC_1_2) + $signed(_zz_io_outputC_1));
  assign _zz__zz_io_outputC_1_2 = {{10{_zz_io_outputC[15]}}, _zz_io_outputC};
  assign io_outputA = io_inputA_regNext;
  assign io_outputB = io_inputB_regNext;
  assign _zz_io_outputC = ($signed(io_inputA) * $signed(io_inputB));
  assign io_outputC = _zz_io_outputC_1;
  always @(posedge clk) begin
    if(reset) begin
      io_inputA_regNext <= 8'h0;
      io_inputB_regNext <= 8'h0;
      _zz_io_outputC_1 <= 26'h0;
    end else begin
      io_inputA_regNext <= io_inputA;
      io_inputB_regNext <= io_inputB;
      _zz_io_outputC_1 <= (io_resetPartialC ? _zz__zz_io_outputC_1 : _zz__zz_io_outputC_1_1);
    end
  end


endmodule
