// Generator : SpinalHDL v1.12.3    git head : 591e64062329e5e2e2b81f4d52422948053edb97
// Component : SInt_ReuseB_SystolicArray_16x16
// Git hash  : c899c5c2103f8885866e344829b479f536941da5

`timescale 1ns/1ps

module SInt_ReuseB_SystolicArray_16x16 (
  input  wire [7:0]    io_inputA_0,
  input  wire [7:0]    io_inputA_1,
  input  wire [7:0]    io_inputA_2,
  input  wire [7:0]    io_inputA_3,
  input  wire [7:0]    io_inputA_4,
  input  wire [7:0]    io_inputA_5,
  input  wire [7:0]    io_inputA_6,
  input  wire [7:0]    io_inputA_7,
  input  wire [7:0]    io_inputA_8,
  input  wire [7:0]    io_inputA_9,
  input  wire [7:0]    io_inputA_10,
  input  wire [7:0]    io_inputA_11,
  input  wire [7:0]    io_inputA_12,
  input  wire [7:0]    io_inputA_13,
  input  wire [7:0]    io_inputA_14,
  input  wire [7:0]    io_inputA_15,
  input  wire [7:0]    io_inputB_0,
  input  wire [7:0]    io_inputB_1,
  input  wire [7:0]    io_inputB_2,
  input  wire [7:0]    io_inputB_3,
  input  wire [7:0]    io_inputB_4,
  input  wire [7:0]    io_inputB_5,
  input  wire [7:0]    io_inputB_6,
  input  wire [7:0]    io_inputB_7,
  input  wire [7:0]    io_inputB_8,
  input  wire [7:0]    io_inputB_9,
  input  wire [7:0]    io_inputB_10,
  input  wire [7:0]    io_inputB_11,
  input  wire [7:0]    io_inputB_12,
  input  wire [7:0]    io_inputB_13,
  input  wire [7:0]    io_inputB_14,
  input  wire [7:0]    io_inputB_15,
  input  wire          io_inputCaptureEnableB_0_0,
  input  wire          io_inputCaptureEnableB_0_1,
  input  wire          io_inputCaptureEnableB_0_2,
  input  wire          io_inputCaptureEnableB_0_3,
  input  wire          io_inputCaptureEnableB_0_4,
  input  wire          io_inputCaptureEnableB_0_5,
  input  wire          io_inputCaptureEnableB_0_6,
  input  wire          io_inputCaptureEnableB_0_7,
  input  wire          io_inputCaptureEnableB_0_8,
  input  wire          io_inputCaptureEnableB_0_9,
  input  wire          io_inputCaptureEnableB_0_10,
  input  wire          io_inputCaptureEnableB_0_11,
  input  wire          io_inputCaptureEnableB_0_12,
  input  wire          io_inputCaptureEnableB_0_13,
  input  wire          io_inputCaptureEnableB_0_14,
  input  wire          io_inputCaptureEnableB_0_15,
  input  wire          io_inputCaptureEnableB_1_0,
  input  wire          io_inputCaptureEnableB_1_1,
  input  wire          io_inputCaptureEnableB_1_2,
  input  wire          io_inputCaptureEnableB_1_3,
  input  wire          io_inputCaptureEnableB_1_4,
  input  wire          io_inputCaptureEnableB_1_5,
  input  wire          io_inputCaptureEnableB_1_6,
  input  wire          io_inputCaptureEnableB_1_7,
  input  wire          io_inputCaptureEnableB_1_8,
  input  wire          io_inputCaptureEnableB_1_9,
  input  wire          io_inputCaptureEnableB_1_10,
  input  wire          io_inputCaptureEnableB_1_11,
  input  wire          io_inputCaptureEnableB_1_12,
  input  wire          io_inputCaptureEnableB_1_13,
  input  wire          io_inputCaptureEnableB_1_14,
  input  wire          io_inputCaptureEnableB_1_15,
  input  wire          io_inputCaptureEnableB_2_0,
  input  wire          io_inputCaptureEnableB_2_1,
  input  wire          io_inputCaptureEnableB_2_2,
  input  wire          io_inputCaptureEnableB_2_3,
  input  wire          io_inputCaptureEnableB_2_4,
  input  wire          io_inputCaptureEnableB_2_5,
  input  wire          io_inputCaptureEnableB_2_6,
  input  wire          io_inputCaptureEnableB_2_7,
  input  wire          io_inputCaptureEnableB_2_8,
  input  wire          io_inputCaptureEnableB_2_9,
  input  wire          io_inputCaptureEnableB_2_10,
  input  wire          io_inputCaptureEnableB_2_11,
  input  wire          io_inputCaptureEnableB_2_12,
  input  wire          io_inputCaptureEnableB_2_13,
  input  wire          io_inputCaptureEnableB_2_14,
  input  wire          io_inputCaptureEnableB_2_15,
  input  wire          io_inputCaptureEnableB_3_0,
  input  wire          io_inputCaptureEnableB_3_1,
  input  wire          io_inputCaptureEnableB_3_2,
  input  wire          io_inputCaptureEnableB_3_3,
  input  wire          io_inputCaptureEnableB_3_4,
  input  wire          io_inputCaptureEnableB_3_5,
  input  wire          io_inputCaptureEnableB_3_6,
  input  wire          io_inputCaptureEnableB_3_7,
  input  wire          io_inputCaptureEnableB_3_8,
  input  wire          io_inputCaptureEnableB_3_9,
  input  wire          io_inputCaptureEnableB_3_10,
  input  wire          io_inputCaptureEnableB_3_11,
  input  wire          io_inputCaptureEnableB_3_12,
  input  wire          io_inputCaptureEnableB_3_13,
  input  wire          io_inputCaptureEnableB_3_14,
  input  wire          io_inputCaptureEnableB_3_15,
  input  wire          io_inputCaptureEnableB_4_0,
  input  wire          io_inputCaptureEnableB_4_1,
  input  wire          io_inputCaptureEnableB_4_2,
  input  wire          io_inputCaptureEnableB_4_3,
  input  wire          io_inputCaptureEnableB_4_4,
  input  wire          io_inputCaptureEnableB_4_5,
  input  wire          io_inputCaptureEnableB_4_6,
  input  wire          io_inputCaptureEnableB_4_7,
  input  wire          io_inputCaptureEnableB_4_8,
  input  wire          io_inputCaptureEnableB_4_9,
  input  wire          io_inputCaptureEnableB_4_10,
  input  wire          io_inputCaptureEnableB_4_11,
  input  wire          io_inputCaptureEnableB_4_12,
  input  wire          io_inputCaptureEnableB_4_13,
  input  wire          io_inputCaptureEnableB_4_14,
  input  wire          io_inputCaptureEnableB_4_15,
  input  wire          io_inputCaptureEnableB_5_0,
  input  wire          io_inputCaptureEnableB_5_1,
  input  wire          io_inputCaptureEnableB_5_2,
  input  wire          io_inputCaptureEnableB_5_3,
  input  wire          io_inputCaptureEnableB_5_4,
  input  wire          io_inputCaptureEnableB_5_5,
  input  wire          io_inputCaptureEnableB_5_6,
  input  wire          io_inputCaptureEnableB_5_7,
  input  wire          io_inputCaptureEnableB_5_8,
  input  wire          io_inputCaptureEnableB_5_9,
  input  wire          io_inputCaptureEnableB_5_10,
  input  wire          io_inputCaptureEnableB_5_11,
  input  wire          io_inputCaptureEnableB_5_12,
  input  wire          io_inputCaptureEnableB_5_13,
  input  wire          io_inputCaptureEnableB_5_14,
  input  wire          io_inputCaptureEnableB_5_15,
  input  wire          io_inputCaptureEnableB_6_0,
  input  wire          io_inputCaptureEnableB_6_1,
  input  wire          io_inputCaptureEnableB_6_2,
  input  wire          io_inputCaptureEnableB_6_3,
  input  wire          io_inputCaptureEnableB_6_4,
  input  wire          io_inputCaptureEnableB_6_5,
  input  wire          io_inputCaptureEnableB_6_6,
  input  wire          io_inputCaptureEnableB_6_7,
  input  wire          io_inputCaptureEnableB_6_8,
  input  wire          io_inputCaptureEnableB_6_9,
  input  wire          io_inputCaptureEnableB_6_10,
  input  wire          io_inputCaptureEnableB_6_11,
  input  wire          io_inputCaptureEnableB_6_12,
  input  wire          io_inputCaptureEnableB_6_13,
  input  wire          io_inputCaptureEnableB_6_14,
  input  wire          io_inputCaptureEnableB_6_15,
  input  wire          io_inputCaptureEnableB_7_0,
  input  wire          io_inputCaptureEnableB_7_1,
  input  wire          io_inputCaptureEnableB_7_2,
  input  wire          io_inputCaptureEnableB_7_3,
  input  wire          io_inputCaptureEnableB_7_4,
  input  wire          io_inputCaptureEnableB_7_5,
  input  wire          io_inputCaptureEnableB_7_6,
  input  wire          io_inputCaptureEnableB_7_7,
  input  wire          io_inputCaptureEnableB_7_8,
  input  wire          io_inputCaptureEnableB_7_9,
  input  wire          io_inputCaptureEnableB_7_10,
  input  wire          io_inputCaptureEnableB_7_11,
  input  wire          io_inputCaptureEnableB_7_12,
  input  wire          io_inputCaptureEnableB_7_13,
  input  wire          io_inputCaptureEnableB_7_14,
  input  wire          io_inputCaptureEnableB_7_15,
  input  wire          io_inputCaptureEnableB_8_0,
  input  wire          io_inputCaptureEnableB_8_1,
  input  wire          io_inputCaptureEnableB_8_2,
  input  wire          io_inputCaptureEnableB_8_3,
  input  wire          io_inputCaptureEnableB_8_4,
  input  wire          io_inputCaptureEnableB_8_5,
  input  wire          io_inputCaptureEnableB_8_6,
  input  wire          io_inputCaptureEnableB_8_7,
  input  wire          io_inputCaptureEnableB_8_8,
  input  wire          io_inputCaptureEnableB_8_9,
  input  wire          io_inputCaptureEnableB_8_10,
  input  wire          io_inputCaptureEnableB_8_11,
  input  wire          io_inputCaptureEnableB_8_12,
  input  wire          io_inputCaptureEnableB_8_13,
  input  wire          io_inputCaptureEnableB_8_14,
  input  wire          io_inputCaptureEnableB_8_15,
  input  wire          io_inputCaptureEnableB_9_0,
  input  wire          io_inputCaptureEnableB_9_1,
  input  wire          io_inputCaptureEnableB_9_2,
  input  wire          io_inputCaptureEnableB_9_3,
  input  wire          io_inputCaptureEnableB_9_4,
  input  wire          io_inputCaptureEnableB_9_5,
  input  wire          io_inputCaptureEnableB_9_6,
  input  wire          io_inputCaptureEnableB_9_7,
  input  wire          io_inputCaptureEnableB_9_8,
  input  wire          io_inputCaptureEnableB_9_9,
  input  wire          io_inputCaptureEnableB_9_10,
  input  wire          io_inputCaptureEnableB_9_11,
  input  wire          io_inputCaptureEnableB_9_12,
  input  wire          io_inputCaptureEnableB_9_13,
  input  wire          io_inputCaptureEnableB_9_14,
  input  wire          io_inputCaptureEnableB_9_15,
  input  wire          io_inputCaptureEnableB_10_0,
  input  wire          io_inputCaptureEnableB_10_1,
  input  wire          io_inputCaptureEnableB_10_2,
  input  wire          io_inputCaptureEnableB_10_3,
  input  wire          io_inputCaptureEnableB_10_4,
  input  wire          io_inputCaptureEnableB_10_5,
  input  wire          io_inputCaptureEnableB_10_6,
  input  wire          io_inputCaptureEnableB_10_7,
  input  wire          io_inputCaptureEnableB_10_8,
  input  wire          io_inputCaptureEnableB_10_9,
  input  wire          io_inputCaptureEnableB_10_10,
  input  wire          io_inputCaptureEnableB_10_11,
  input  wire          io_inputCaptureEnableB_10_12,
  input  wire          io_inputCaptureEnableB_10_13,
  input  wire          io_inputCaptureEnableB_10_14,
  input  wire          io_inputCaptureEnableB_10_15,
  input  wire          io_inputCaptureEnableB_11_0,
  input  wire          io_inputCaptureEnableB_11_1,
  input  wire          io_inputCaptureEnableB_11_2,
  input  wire          io_inputCaptureEnableB_11_3,
  input  wire          io_inputCaptureEnableB_11_4,
  input  wire          io_inputCaptureEnableB_11_5,
  input  wire          io_inputCaptureEnableB_11_6,
  input  wire          io_inputCaptureEnableB_11_7,
  input  wire          io_inputCaptureEnableB_11_8,
  input  wire          io_inputCaptureEnableB_11_9,
  input  wire          io_inputCaptureEnableB_11_10,
  input  wire          io_inputCaptureEnableB_11_11,
  input  wire          io_inputCaptureEnableB_11_12,
  input  wire          io_inputCaptureEnableB_11_13,
  input  wire          io_inputCaptureEnableB_11_14,
  input  wire          io_inputCaptureEnableB_11_15,
  input  wire          io_inputCaptureEnableB_12_0,
  input  wire          io_inputCaptureEnableB_12_1,
  input  wire          io_inputCaptureEnableB_12_2,
  input  wire          io_inputCaptureEnableB_12_3,
  input  wire          io_inputCaptureEnableB_12_4,
  input  wire          io_inputCaptureEnableB_12_5,
  input  wire          io_inputCaptureEnableB_12_6,
  input  wire          io_inputCaptureEnableB_12_7,
  input  wire          io_inputCaptureEnableB_12_8,
  input  wire          io_inputCaptureEnableB_12_9,
  input  wire          io_inputCaptureEnableB_12_10,
  input  wire          io_inputCaptureEnableB_12_11,
  input  wire          io_inputCaptureEnableB_12_12,
  input  wire          io_inputCaptureEnableB_12_13,
  input  wire          io_inputCaptureEnableB_12_14,
  input  wire          io_inputCaptureEnableB_12_15,
  input  wire          io_inputCaptureEnableB_13_0,
  input  wire          io_inputCaptureEnableB_13_1,
  input  wire          io_inputCaptureEnableB_13_2,
  input  wire          io_inputCaptureEnableB_13_3,
  input  wire          io_inputCaptureEnableB_13_4,
  input  wire          io_inputCaptureEnableB_13_5,
  input  wire          io_inputCaptureEnableB_13_6,
  input  wire          io_inputCaptureEnableB_13_7,
  input  wire          io_inputCaptureEnableB_13_8,
  input  wire          io_inputCaptureEnableB_13_9,
  input  wire          io_inputCaptureEnableB_13_10,
  input  wire          io_inputCaptureEnableB_13_11,
  input  wire          io_inputCaptureEnableB_13_12,
  input  wire          io_inputCaptureEnableB_13_13,
  input  wire          io_inputCaptureEnableB_13_14,
  input  wire          io_inputCaptureEnableB_13_15,
  input  wire          io_inputCaptureEnableB_14_0,
  input  wire          io_inputCaptureEnableB_14_1,
  input  wire          io_inputCaptureEnableB_14_2,
  input  wire          io_inputCaptureEnableB_14_3,
  input  wire          io_inputCaptureEnableB_14_4,
  input  wire          io_inputCaptureEnableB_14_5,
  input  wire          io_inputCaptureEnableB_14_6,
  input  wire          io_inputCaptureEnableB_14_7,
  input  wire          io_inputCaptureEnableB_14_8,
  input  wire          io_inputCaptureEnableB_14_9,
  input  wire          io_inputCaptureEnableB_14_10,
  input  wire          io_inputCaptureEnableB_14_11,
  input  wire          io_inputCaptureEnableB_14_12,
  input  wire          io_inputCaptureEnableB_14_13,
  input  wire          io_inputCaptureEnableB_14_14,
  input  wire          io_inputCaptureEnableB_14_15,
  input  wire          io_inputCaptureEnableB_15_0,
  input  wire          io_inputCaptureEnableB_15_1,
  input  wire          io_inputCaptureEnableB_15_2,
  input  wire          io_inputCaptureEnableB_15_3,
  input  wire          io_inputCaptureEnableB_15_4,
  input  wire          io_inputCaptureEnableB_15_5,
  input  wire          io_inputCaptureEnableB_15_6,
  input  wire          io_inputCaptureEnableB_15_7,
  input  wire          io_inputCaptureEnableB_15_8,
  input  wire          io_inputCaptureEnableB_15_9,
  input  wire          io_inputCaptureEnableB_15_10,
  input  wire          io_inputCaptureEnableB_15_11,
  input  wire          io_inputCaptureEnableB_15_12,
  input  wire          io_inputCaptureEnableB_15_13,
  input  wire          io_inputCaptureEnableB_15_14,
  input  wire          io_inputCaptureEnableB_15_15,
  output wire [19:0]   io_outputC_0,
  output wire [19:0]   io_outputC_1,
  output wire [19:0]   io_outputC_2,
  output wire [19:0]   io_outputC_3,
  output wire [19:0]   io_outputC_4,
  output wire [19:0]   io_outputC_5,
  output wire [19:0]   io_outputC_6,
  output wire [19:0]   io_outputC_7,
  output wire [19:0]   io_outputC_8,
  output wire [19:0]   io_outputC_9,
  output wire [19:0]   io_outputC_10,
  output wire [19:0]   io_outputC_11,
  output wire [19:0]   io_outputC_12,
  output wire [19:0]   io_outputC_13,
  output wire [19:0]   io_outputC_14,
  output wire [19:0]   io_outputC_15,
  input  wire          clk,
  input  wire          reset
);
//#region Internal Wires/Regs
  wire       [7:0]    pes_0_0_io_outputA;
  wire       [7:0]    pes_0_0_io_outputB;
  wire       [15:0]   pes_0_0_io_outputC;
  wire       [7:0]    pes_0_1_io_outputA;
  wire       [7:0]    pes_0_1_io_outputB;
  wire       [15:0]   pes_0_1_io_outputC;
  wire       [7:0]    pes_0_2_io_outputA;
  wire       [7:0]    pes_0_2_io_outputB;
  wire       [15:0]   pes_0_2_io_outputC;
  wire       [7:0]    pes_0_3_io_outputA;
  wire       [7:0]    pes_0_3_io_outputB;
  wire       [15:0]   pes_0_3_io_outputC;
  wire       [7:0]    pes_0_4_io_outputA;
  wire       [7:0]    pes_0_4_io_outputB;
  wire       [15:0]   pes_0_4_io_outputC;
  wire       [7:0]    pes_0_5_io_outputA;
  wire       [7:0]    pes_0_5_io_outputB;
  wire       [15:0]   pes_0_5_io_outputC;
  wire       [7:0]    pes_0_6_io_outputA;
  wire       [7:0]    pes_0_6_io_outputB;
  wire       [15:0]   pes_0_6_io_outputC;
  wire       [7:0]    pes_0_7_io_outputA;
  wire       [7:0]    pes_0_7_io_outputB;
  wire       [15:0]   pes_0_7_io_outputC;
  wire       [7:0]    pes_0_8_io_outputA;
  wire       [7:0]    pes_0_8_io_outputB;
  wire       [15:0]   pes_0_8_io_outputC;
  wire       [7:0]    pes_0_9_io_outputA;
  wire       [7:0]    pes_0_9_io_outputB;
  wire       [15:0]   pes_0_9_io_outputC;
  wire       [7:0]    pes_0_10_io_outputA;
  wire       [7:0]    pes_0_10_io_outputB;
  wire       [15:0]   pes_0_10_io_outputC;
  wire       [7:0]    pes_0_11_io_outputA;
  wire       [7:0]    pes_0_11_io_outputB;
  wire       [15:0]   pes_0_11_io_outputC;
  wire       [7:0]    pes_0_12_io_outputA;
  wire       [7:0]    pes_0_12_io_outputB;
  wire       [15:0]   pes_0_12_io_outputC;
  wire       [7:0]    pes_0_13_io_outputA;
  wire       [7:0]    pes_0_13_io_outputB;
  wire       [15:0]   pes_0_13_io_outputC;
  wire       [7:0]    pes_0_14_io_outputA;
  wire       [7:0]    pes_0_14_io_outputB;
  wire       [15:0]   pes_0_14_io_outputC;
  wire       [7:0]    pes_0_15_io_outputB;
  wire       [15:0]   pes_0_15_io_outputC;
  wire       [7:0]    pes_1_0_io_outputA;
  wire       [7:0]    pes_1_0_io_outputB;
  wire       [16:0]   pes_1_0_io_outputC;
  wire       [7:0]    pes_1_1_io_outputA;
  wire       [7:0]    pes_1_1_io_outputB;
  wire       [16:0]   pes_1_1_io_outputC;
  wire       [7:0]    pes_1_2_io_outputA;
  wire       [7:0]    pes_1_2_io_outputB;
  wire       [16:0]   pes_1_2_io_outputC;
  wire       [7:0]    pes_1_3_io_outputA;
  wire       [7:0]    pes_1_3_io_outputB;
  wire       [16:0]   pes_1_3_io_outputC;
  wire       [7:0]    pes_1_4_io_outputA;
  wire       [7:0]    pes_1_4_io_outputB;
  wire       [16:0]   pes_1_4_io_outputC;
  wire       [7:0]    pes_1_5_io_outputA;
  wire       [7:0]    pes_1_5_io_outputB;
  wire       [16:0]   pes_1_5_io_outputC;
  wire       [7:0]    pes_1_6_io_outputA;
  wire       [7:0]    pes_1_6_io_outputB;
  wire       [16:0]   pes_1_6_io_outputC;
  wire       [7:0]    pes_1_7_io_outputA;
  wire       [7:0]    pes_1_7_io_outputB;
  wire       [16:0]   pes_1_7_io_outputC;
  wire       [7:0]    pes_1_8_io_outputA;
  wire       [7:0]    pes_1_8_io_outputB;
  wire       [16:0]   pes_1_8_io_outputC;
  wire       [7:0]    pes_1_9_io_outputA;
  wire       [7:0]    pes_1_9_io_outputB;
  wire       [16:0]   pes_1_9_io_outputC;
  wire       [7:0]    pes_1_10_io_outputA;
  wire       [7:0]    pes_1_10_io_outputB;
  wire       [16:0]   pes_1_10_io_outputC;
  wire       [7:0]    pes_1_11_io_outputA;
  wire       [7:0]    pes_1_11_io_outputB;
  wire       [16:0]   pes_1_11_io_outputC;
  wire       [7:0]    pes_1_12_io_outputA;
  wire       [7:0]    pes_1_12_io_outputB;
  wire       [16:0]   pes_1_12_io_outputC;
  wire       [7:0]    pes_1_13_io_outputA;
  wire       [7:0]    pes_1_13_io_outputB;
  wire       [16:0]   pes_1_13_io_outputC;
  wire       [7:0]    pes_1_14_io_outputA;
  wire       [7:0]    pes_1_14_io_outputB;
  wire       [16:0]   pes_1_14_io_outputC;
  wire       [7:0]    pes_1_15_io_outputB;
  wire       [16:0]   pes_1_15_io_outputC;
  wire       [7:0]    pes_2_0_io_outputA;
  wire       [7:0]    pes_2_0_io_outputB;
  wire       [17:0]   pes_2_0_io_outputC;
  wire       [7:0]    pes_2_1_io_outputA;
  wire       [7:0]    pes_2_1_io_outputB;
  wire       [17:0]   pes_2_1_io_outputC;
  wire       [7:0]    pes_2_2_io_outputA;
  wire       [7:0]    pes_2_2_io_outputB;
  wire       [17:0]   pes_2_2_io_outputC;
  wire       [7:0]    pes_2_3_io_outputA;
  wire       [7:0]    pes_2_3_io_outputB;
  wire       [17:0]   pes_2_3_io_outputC;
  wire       [7:0]    pes_2_4_io_outputA;
  wire       [7:0]    pes_2_4_io_outputB;
  wire       [17:0]   pes_2_4_io_outputC;
  wire       [7:0]    pes_2_5_io_outputA;
  wire       [7:0]    pes_2_5_io_outputB;
  wire       [17:0]   pes_2_5_io_outputC;
  wire       [7:0]    pes_2_6_io_outputA;
  wire       [7:0]    pes_2_6_io_outputB;
  wire       [17:0]   pes_2_6_io_outputC;
  wire       [7:0]    pes_2_7_io_outputA;
  wire       [7:0]    pes_2_7_io_outputB;
  wire       [17:0]   pes_2_7_io_outputC;
  wire       [7:0]    pes_2_8_io_outputA;
  wire       [7:0]    pes_2_8_io_outputB;
  wire       [17:0]   pes_2_8_io_outputC;
  wire       [7:0]    pes_2_9_io_outputA;
  wire       [7:0]    pes_2_9_io_outputB;
  wire       [17:0]   pes_2_9_io_outputC;
  wire       [7:0]    pes_2_10_io_outputA;
  wire       [7:0]    pes_2_10_io_outputB;
  wire       [17:0]   pes_2_10_io_outputC;
  wire       [7:0]    pes_2_11_io_outputA;
  wire       [7:0]    pes_2_11_io_outputB;
  wire       [17:0]   pes_2_11_io_outputC;
  wire       [7:0]    pes_2_12_io_outputA;
  wire       [7:0]    pes_2_12_io_outputB;
  wire       [17:0]   pes_2_12_io_outputC;
  wire       [7:0]    pes_2_13_io_outputA;
  wire       [7:0]    pes_2_13_io_outputB;
  wire       [17:0]   pes_2_13_io_outputC;
  wire       [7:0]    pes_2_14_io_outputA;
  wire       [7:0]    pes_2_14_io_outputB;
  wire       [17:0]   pes_2_14_io_outputC;
  wire       [7:0]    pes_2_15_io_outputB;
  wire       [17:0]   pes_2_15_io_outputC;
  wire       [7:0]    pes_3_0_io_outputA;
  wire       [7:0]    pes_3_0_io_outputB;
  wire       [17:0]   pes_3_0_io_outputC;
  wire       [7:0]    pes_3_1_io_outputA;
  wire       [7:0]    pes_3_1_io_outputB;
  wire       [17:0]   pes_3_1_io_outputC;
  wire       [7:0]    pes_3_2_io_outputA;
  wire       [7:0]    pes_3_2_io_outputB;
  wire       [17:0]   pes_3_2_io_outputC;
  wire       [7:0]    pes_3_3_io_outputA;
  wire       [7:0]    pes_3_3_io_outputB;
  wire       [17:0]   pes_3_3_io_outputC;
  wire       [7:0]    pes_3_4_io_outputA;
  wire       [7:0]    pes_3_4_io_outputB;
  wire       [17:0]   pes_3_4_io_outputC;
  wire       [7:0]    pes_3_5_io_outputA;
  wire       [7:0]    pes_3_5_io_outputB;
  wire       [17:0]   pes_3_5_io_outputC;
  wire       [7:0]    pes_3_6_io_outputA;
  wire       [7:0]    pes_3_6_io_outputB;
  wire       [17:0]   pes_3_6_io_outputC;
  wire       [7:0]    pes_3_7_io_outputA;
  wire       [7:0]    pes_3_7_io_outputB;
  wire       [17:0]   pes_3_7_io_outputC;
  wire       [7:0]    pes_3_8_io_outputA;
  wire       [7:0]    pes_3_8_io_outputB;
  wire       [17:0]   pes_3_8_io_outputC;
  wire       [7:0]    pes_3_9_io_outputA;
  wire       [7:0]    pes_3_9_io_outputB;
  wire       [17:0]   pes_3_9_io_outputC;
  wire       [7:0]    pes_3_10_io_outputA;
  wire       [7:0]    pes_3_10_io_outputB;
  wire       [17:0]   pes_3_10_io_outputC;
  wire       [7:0]    pes_3_11_io_outputA;
  wire       [7:0]    pes_3_11_io_outputB;
  wire       [17:0]   pes_3_11_io_outputC;
  wire       [7:0]    pes_3_12_io_outputA;
  wire       [7:0]    pes_3_12_io_outputB;
  wire       [17:0]   pes_3_12_io_outputC;
  wire       [7:0]    pes_3_13_io_outputA;
  wire       [7:0]    pes_3_13_io_outputB;
  wire       [17:0]   pes_3_13_io_outputC;
  wire       [7:0]    pes_3_14_io_outputA;
  wire       [7:0]    pes_3_14_io_outputB;
  wire       [17:0]   pes_3_14_io_outputC;
  wire       [7:0]    pes_3_15_io_outputB;
  wire       [17:0]   pes_3_15_io_outputC;
  wire       [7:0]    pes_4_0_io_outputA;
  wire       [7:0]    pes_4_0_io_outputB;
  wire       [18:0]   pes_4_0_io_outputC;
  wire       [7:0]    pes_4_1_io_outputA;
  wire       [7:0]    pes_4_1_io_outputB;
  wire       [18:0]   pes_4_1_io_outputC;
  wire       [7:0]    pes_4_2_io_outputA;
  wire       [7:0]    pes_4_2_io_outputB;
  wire       [18:0]   pes_4_2_io_outputC;
  wire       [7:0]    pes_4_3_io_outputA;
  wire       [7:0]    pes_4_3_io_outputB;
  wire       [18:0]   pes_4_3_io_outputC;
  wire       [7:0]    pes_4_4_io_outputA;
  wire       [7:0]    pes_4_4_io_outputB;
  wire       [18:0]   pes_4_4_io_outputC;
  wire       [7:0]    pes_4_5_io_outputA;
  wire       [7:0]    pes_4_5_io_outputB;
  wire       [18:0]   pes_4_5_io_outputC;
  wire       [7:0]    pes_4_6_io_outputA;
  wire       [7:0]    pes_4_6_io_outputB;
  wire       [18:0]   pes_4_6_io_outputC;
  wire       [7:0]    pes_4_7_io_outputA;
  wire       [7:0]    pes_4_7_io_outputB;
  wire       [18:0]   pes_4_7_io_outputC;
  wire       [7:0]    pes_4_8_io_outputA;
  wire       [7:0]    pes_4_8_io_outputB;
  wire       [18:0]   pes_4_8_io_outputC;
  wire       [7:0]    pes_4_9_io_outputA;
  wire       [7:0]    pes_4_9_io_outputB;
  wire       [18:0]   pes_4_9_io_outputC;
  wire       [7:0]    pes_4_10_io_outputA;
  wire       [7:0]    pes_4_10_io_outputB;
  wire       [18:0]   pes_4_10_io_outputC;
  wire       [7:0]    pes_4_11_io_outputA;
  wire       [7:0]    pes_4_11_io_outputB;
  wire       [18:0]   pes_4_11_io_outputC;
  wire       [7:0]    pes_4_12_io_outputA;
  wire       [7:0]    pes_4_12_io_outputB;
  wire       [18:0]   pes_4_12_io_outputC;
  wire       [7:0]    pes_4_13_io_outputA;
  wire       [7:0]    pes_4_13_io_outputB;
  wire       [18:0]   pes_4_13_io_outputC;
  wire       [7:0]    pes_4_14_io_outputA;
  wire       [7:0]    pes_4_14_io_outputB;
  wire       [18:0]   pes_4_14_io_outputC;
  wire       [7:0]    pes_4_15_io_outputB;
  wire       [18:0]   pes_4_15_io_outputC;
  wire       [7:0]    pes_5_0_io_outputA;
  wire       [7:0]    pes_5_0_io_outputB;
  wire       [18:0]   pes_5_0_io_outputC;
  wire       [7:0]    pes_5_1_io_outputA;
  wire       [7:0]    pes_5_1_io_outputB;
  wire       [18:0]   pes_5_1_io_outputC;
  wire       [7:0]    pes_5_2_io_outputA;
  wire       [7:0]    pes_5_2_io_outputB;
  wire       [18:0]   pes_5_2_io_outputC;
  wire       [7:0]    pes_5_3_io_outputA;
  wire       [7:0]    pes_5_3_io_outputB;
  wire       [18:0]   pes_5_3_io_outputC;
  wire       [7:0]    pes_5_4_io_outputA;
  wire       [7:0]    pes_5_4_io_outputB;
  wire       [18:0]   pes_5_4_io_outputC;
  wire       [7:0]    pes_5_5_io_outputA;
  wire       [7:0]    pes_5_5_io_outputB;
  wire       [18:0]   pes_5_5_io_outputC;
  wire       [7:0]    pes_5_6_io_outputA;
  wire       [7:0]    pes_5_6_io_outputB;
  wire       [18:0]   pes_5_6_io_outputC;
  wire       [7:0]    pes_5_7_io_outputA;
  wire       [7:0]    pes_5_7_io_outputB;
  wire       [18:0]   pes_5_7_io_outputC;
  wire       [7:0]    pes_5_8_io_outputA;
  wire       [7:0]    pes_5_8_io_outputB;
  wire       [18:0]   pes_5_8_io_outputC;
  wire       [7:0]    pes_5_9_io_outputA;
  wire       [7:0]    pes_5_9_io_outputB;
  wire       [18:0]   pes_5_9_io_outputC;
  wire       [7:0]    pes_5_10_io_outputA;
  wire       [7:0]    pes_5_10_io_outputB;
  wire       [18:0]   pes_5_10_io_outputC;
  wire       [7:0]    pes_5_11_io_outputA;
  wire       [7:0]    pes_5_11_io_outputB;
  wire       [18:0]   pes_5_11_io_outputC;
  wire       [7:0]    pes_5_12_io_outputA;
  wire       [7:0]    pes_5_12_io_outputB;
  wire       [18:0]   pes_5_12_io_outputC;
  wire       [7:0]    pes_5_13_io_outputA;
  wire       [7:0]    pes_5_13_io_outputB;
  wire       [18:0]   pes_5_13_io_outputC;
  wire       [7:0]    pes_5_14_io_outputA;
  wire       [7:0]    pes_5_14_io_outputB;
  wire       [18:0]   pes_5_14_io_outputC;
  wire       [7:0]    pes_5_15_io_outputB;
  wire       [18:0]   pes_5_15_io_outputC;
  wire       [7:0]    pes_6_0_io_outputA;
  wire       [7:0]    pes_6_0_io_outputB;
  wire       [18:0]   pes_6_0_io_outputC;
  wire       [7:0]    pes_6_1_io_outputA;
  wire       [7:0]    pes_6_1_io_outputB;
  wire       [18:0]   pes_6_1_io_outputC;
  wire       [7:0]    pes_6_2_io_outputA;
  wire       [7:0]    pes_6_2_io_outputB;
  wire       [18:0]   pes_6_2_io_outputC;
  wire       [7:0]    pes_6_3_io_outputA;
  wire       [7:0]    pes_6_3_io_outputB;
  wire       [18:0]   pes_6_3_io_outputC;
  wire       [7:0]    pes_6_4_io_outputA;
  wire       [7:0]    pes_6_4_io_outputB;
  wire       [18:0]   pes_6_4_io_outputC;
  wire       [7:0]    pes_6_5_io_outputA;
  wire       [7:0]    pes_6_5_io_outputB;
  wire       [18:0]   pes_6_5_io_outputC;
  wire       [7:0]    pes_6_6_io_outputA;
  wire       [7:0]    pes_6_6_io_outputB;
  wire       [18:0]   pes_6_6_io_outputC;
  wire       [7:0]    pes_6_7_io_outputA;
  wire       [7:0]    pes_6_7_io_outputB;
  wire       [18:0]   pes_6_7_io_outputC;
  wire       [7:0]    pes_6_8_io_outputA;
  wire       [7:0]    pes_6_8_io_outputB;
  wire       [18:0]   pes_6_8_io_outputC;
  wire       [7:0]    pes_6_9_io_outputA;
  wire       [7:0]    pes_6_9_io_outputB;
  wire       [18:0]   pes_6_9_io_outputC;
  wire       [7:0]    pes_6_10_io_outputA;
  wire       [7:0]    pes_6_10_io_outputB;
  wire       [18:0]   pes_6_10_io_outputC;
  wire       [7:0]    pes_6_11_io_outputA;
  wire       [7:0]    pes_6_11_io_outputB;
  wire       [18:0]   pes_6_11_io_outputC;
  wire       [7:0]    pes_6_12_io_outputA;
  wire       [7:0]    pes_6_12_io_outputB;
  wire       [18:0]   pes_6_12_io_outputC;
  wire       [7:0]    pes_6_13_io_outputA;
  wire       [7:0]    pes_6_13_io_outputB;
  wire       [18:0]   pes_6_13_io_outputC;
  wire       [7:0]    pes_6_14_io_outputA;
  wire       [7:0]    pes_6_14_io_outputB;
  wire       [18:0]   pes_6_14_io_outputC;
  wire       [7:0]    pes_6_15_io_outputB;
  wire       [18:0]   pes_6_15_io_outputC;
  wire       [7:0]    pes_7_0_io_outputA;
  wire       [7:0]    pes_7_0_io_outputB;
  wire       [18:0]   pes_7_0_io_outputC;
  wire       [7:0]    pes_7_1_io_outputA;
  wire       [7:0]    pes_7_1_io_outputB;
  wire       [18:0]   pes_7_1_io_outputC;
  wire       [7:0]    pes_7_2_io_outputA;
  wire       [7:0]    pes_7_2_io_outputB;
  wire       [18:0]   pes_7_2_io_outputC;
  wire       [7:0]    pes_7_3_io_outputA;
  wire       [7:0]    pes_7_3_io_outputB;
  wire       [18:0]   pes_7_3_io_outputC;
  wire       [7:0]    pes_7_4_io_outputA;
  wire       [7:0]    pes_7_4_io_outputB;
  wire       [18:0]   pes_7_4_io_outputC;
  wire       [7:0]    pes_7_5_io_outputA;
  wire       [7:0]    pes_7_5_io_outputB;
  wire       [18:0]   pes_7_5_io_outputC;
  wire       [7:0]    pes_7_6_io_outputA;
  wire       [7:0]    pes_7_6_io_outputB;
  wire       [18:0]   pes_7_6_io_outputC;
  wire       [7:0]    pes_7_7_io_outputA;
  wire       [7:0]    pes_7_7_io_outputB;
  wire       [18:0]   pes_7_7_io_outputC;
  wire       [7:0]    pes_7_8_io_outputA;
  wire       [7:0]    pes_7_8_io_outputB;
  wire       [18:0]   pes_7_8_io_outputC;
  wire       [7:0]    pes_7_9_io_outputA;
  wire       [7:0]    pes_7_9_io_outputB;
  wire       [18:0]   pes_7_9_io_outputC;
  wire       [7:0]    pes_7_10_io_outputA;
  wire       [7:0]    pes_7_10_io_outputB;
  wire       [18:0]   pes_7_10_io_outputC;
  wire       [7:0]    pes_7_11_io_outputA;
  wire       [7:0]    pes_7_11_io_outputB;
  wire       [18:0]   pes_7_11_io_outputC;
  wire       [7:0]    pes_7_12_io_outputA;
  wire       [7:0]    pes_7_12_io_outputB;
  wire       [18:0]   pes_7_12_io_outputC;
  wire       [7:0]    pes_7_13_io_outputA;
  wire       [7:0]    pes_7_13_io_outputB;
  wire       [18:0]   pes_7_13_io_outputC;
  wire       [7:0]    pes_7_14_io_outputA;
  wire       [7:0]    pes_7_14_io_outputB;
  wire       [18:0]   pes_7_14_io_outputC;
  wire       [7:0]    pes_7_15_io_outputB;
  wire       [18:0]   pes_7_15_io_outputC;
  wire       [7:0]    pes_8_0_io_outputA;
  wire       [7:0]    pes_8_0_io_outputB;
  wire       [19:0]   pes_8_0_io_outputC;
  wire       [7:0]    pes_8_1_io_outputA;
  wire       [7:0]    pes_8_1_io_outputB;
  wire       [19:0]   pes_8_1_io_outputC;
  wire       [7:0]    pes_8_2_io_outputA;
  wire       [7:0]    pes_8_2_io_outputB;
  wire       [19:0]   pes_8_2_io_outputC;
  wire       [7:0]    pes_8_3_io_outputA;
  wire       [7:0]    pes_8_3_io_outputB;
  wire       [19:0]   pes_8_3_io_outputC;
  wire       [7:0]    pes_8_4_io_outputA;
  wire       [7:0]    pes_8_4_io_outputB;
  wire       [19:0]   pes_8_4_io_outputC;
  wire       [7:0]    pes_8_5_io_outputA;
  wire       [7:0]    pes_8_5_io_outputB;
  wire       [19:0]   pes_8_5_io_outputC;
  wire       [7:0]    pes_8_6_io_outputA;
  wire       [7:0]    pes_8_6_io_outputB;
  wire       [19:0]   pes_8_6_io_outputC;
  wire       [7:0]    pes_8_7_io_outputA;
  wire       [7:0]    pes_8_7_io_outputB;
  wire       [19:0]   pes_8_7_io_outputC;
  wire       [7:0]    pes_8_8_io_outputA;
  wire       [7:0]    pes_8_8_io_outputB;
  wire       [19:0]   pes_8_8_io_outputC;
  wire       [7:0]    pes_8_9_io_outputA;
  wire       [7:0]    pes_8_9_io_outputB;
  wire       [19:0]   pes_8_9_io_outputC;
  wire       [7:0]    pes_8_10_io_outputA;
  wire       [7:0]    pes_8_10_io_outputB;
  wire       [19:0]   pes_8_10_io_outputC;
  wire       [7:0]    pes_8_11_io_outputA;
  wire       [7:0]    pes_8_11_io_outputB;
  wire       [19:0]   pes_8_11_io_outputC;
  wire       [7:0]    pes_8_12_io_outputA;
  wire       [7:0]    pes_8_12_io_outputB;
  wire       [19:0]   pes_8_12_io_outputC;
  wire       [7:0]    pes_8_13_io_outputA;
  wire       [7:0]    pes_8_13_io_outputB;
  wire       [19:0]   pes_8_13_io_outputC;
  wire       [7:0]    pes_8_14_io_outputA;
  wire       [7:0]    pes_8_14_io_outputB;
  wire       [19:0]   pes_8_14_io_outputC;
  wire       [7:0]    pes_8_15_io_outputB;
  wire       [19:0]   pes_8_15_io_outputC;
  wire       [7:0]    pes_9_0_io_outputA;
  wire       [7:0]    pes_9_0_io_outputB;
  wire       [19:0]   pes_9_0_io_outputC;
  wire       [7:0]    pes_9_1_io_outputA;
  wire       [7:0]    pes_9_1_io_outputB;
  wire       [19:0]   pes_9_1_io_outputC;
  wire       [7:0]    pes_9_2_io_outputA;
  wire       [7:0]    pes_9_2_io_outputB;
  wire       [19:0]   pes_9_2_io_outputC;
  wire       [7:0]    pes_9_3_io_outputA;
  wire       [7:0]    pes_9_3_io_outputB;
  wire       [19:0]   pes_9_3_io_outputC;
  wire       [7:0]    pes_9_4_io_outputA;
  wire       [7:0]    pes_9_4_io_outputB;
  wire       [19:0]   pes_9_4_io_outputC;
  wire       [7:0]    pes_9_5_io_outputA;
  wire       [7:0]    pes_9_5_io_outputB;
  wire       [19:0]   pes_9_5_io_outputC;
  wire       [7:0]    pes_9_6_io_outputA;
  wire       [7:0]    pes_9_6_io_outputB;
  wire       [19:0]   pes_9_6_io_outputC;
  wire       [7:0]    pes_9_7_io_outputA;
  wire       [7:0]    pes_9_7_io_outputB;
  wire       [19:0]   pes_9_7_io_outputC;
  wire       [7:0]    pes_9_8_io_outputA;
  wire       [7:0]    pes_9_8_io_outputB;
  wire       [19:0]   pes_9_8_io_outputC;
  wire       [7:0]    pes_9_9_io_outputA;
  wire       [7:0]    pes_9_9_io_outputB;
  wire       [19:0]   pes_9_9_io_outputC;
  wire       [7:0]    pes_9_10_io_outputA;
  wire       [7:0]    pes_9_10_io_outputB;
  wire       [19:0]   pes_9_10_io_outputC;
  wire       [7:0]    pes_9_11_io_outputA;
  wire       [7:0]    pes_9_11_io_outputB;
  wire       [19:0]   pes_9_11_io_outputC;
  wire       [7:0]    pes_9_12_io_outputA;
  wire       [7:0]    pes_9_12_io_outputB;
  wire       [19:0]   pes_9_12_io_outputC;
  wire       [7:0]    pes_9_13_io_outputA;
  wire       [7:0]    pes_9_13_io_outputB;
  wire       [19:0]   pes_9_13_io_outputC;
  wire       [7:0]    pes_9_14_io_outputA;
  wire       [7:0]    pes_9_14_io_outputB;
  wire       [19:0]   pes_9_14_io_outputC;
  wire       [7:0]    pes_9_15_io_outputB;
  wire       [19:0]   pes_9_15_io_outputC;
  wire       [7:0]    pes_10_0_io_outputA;
  wire       [7:0]    pes_10_0_io_outputB;
  wire       [19:0]   pes_10_0_io_outputC;
  wire       [7:0]    pes_10_1_io_outputA;
  wire       [7:0]    pes_10_1_io_outputB;
  wire       [19:0]   pes_10_1_io_outputC;
  wire       [7:0]    pes_10_2_io_outputA;
  wire       [7:0]    pes_10_2_io_outputB;
  wire       [19:0]   pes_10_2_io_outputC;
  wire       [7:0]    pes_10_3_io_outputA;
  wire       [7:0]    pes_10_3_io_outputB;
  wire       [19:0]   pes_10_3_io_outputC;
  wire       [7:0]    pes_10_4_io_outputA;
  wire       [7:0]    pes_10_4_io_outputB;
  wire       [19:0]   pes_10_4_io_outputC;
  wire       [7:0]    pes_10_5_io_outputA;
  wire       [7:0]    pes_10_5_io_outputB;
  wire       [19:0]   pes_10_5_io_outputC;
  wire       [7:0]    pes_10_6_io_outputA;
  wire       [7:0]    pes_10_6_io_outputB;
  wire       [19:0]   pes_10_6_io_outputC;
  wire       [7:0]    pes_10_7_io_outputA;
  wire       [7:0]    pes_10_7_io_outputB;
  wire       [19:0]   pes_10_7_io_outputC;
  wire       [7:0]    pes_10_8_io_outputA;
  wire       [7:0]    pes_10_8_io_outputB;
  wire       [19:0]   pes_10_8_io_outputC;
  wire       [7:0]    pes_10_9_io_outputA;
  wire       [7:0]    pes_10_9_io_outputB;
  wire       [19:0]   pes_10_9_io_outputC;
  wire       [7:0]    pes_10_10_io_outputA;
  wire       [7:0]    pes_10_10_io_outputB;
  wire       [19:0]   pes_10_10_io_outputC;
  wire       [7:0]    pes_10_11_io_outputA;
  wire       [7:0]    pes_10_11_io_outputB;
  wire       [19:0]   pes_10_11_io_outputC;
  wire       [7:0]    pes_10_12_io_outputA;
  wire       [7:0]    pes_10_12_io_outputB;
  wire       [19:0]   pes_10_12_io_outputC;
  wire       [7:0]    pes_10_13_io_outputA;
  wire       [7:0]    pes_10_13_io_outputB;
  wire       [19:0]   pes_10_13_io_outputC;
  wire       [7:0]    pes_10_14_io_outputA;
  wire       [7:0]    pes_10_14_io_outputB;
  wire       [19:0]   pes_10_14_io_outputC;
  wire       [7:0]    pes_10_15_io_outputB;
  wire       [19:0]   pes_10_15_io_outputC;
  wire       [7:0]    pes_11_0_io_outputA;
  wire       [7:0]    pes_11_0_io_outputB;
  wire       [19:0]   pes_11_0_io_outputC;
  wire       [7:0]    pes_11_1_io_outputA;
  wire       [7:0]    pes_11_1_io_outputB;
  wire       [19:0]   pes_11_1_io_outputC;
  wire       [7:0]    pes_11_2_io_outputA;
  wire       [7:0]    pes_11_2_io_outputB;
  wire       [19:0]   pes_11_2_io_outputC;
  wire       [7:0]    pes_11_3_io_outputA;
  wire       [7:0]    pes_11_3_io_outputB;
  wire       [19:0]   pes_11_3_io_outputC;
  wire       [7:0]    pes_11_4_io_outputA;
  wire       [7:0]    pes_11_4_io_outputB;
  wire       [19:0]   pes_11_4_io_outputC;
  wire       [7:0]    pes_11_5_io_outputA;
  wire       [7:0]    pes_11_5_io_outputB;
  wire       [19:0]   pes_11_5_io_outputC;
  wire       [7:0]    pes_11_6_io_outputA;
  wire       [7:0]    pes_11_6_io_outputB;
  wire       [19:0]   pes_11_6_io_outputC;
  wire       [7:0]    pes_11_7_io_outputA;
  wire       [7:0]    pes_11_7_io_outputB;
  wire       [19:0]   pes_11_7_io_outputC;
  wire       [7:0]    pes_11_8_io_outputA;
  wire       [7:0]    pes_11_8_io_outputB;
  wire       [19:0]   pes_11_8_io_outputC;
  wire       [7:0]    pes_11_9_io_outputA;
  wire       [7:0]    pes_11_9_io_outputB;
  wire       [19:0]   pes_11_9_io_outputC;
  wire       [7:0]    pes_11_10_io_outputA;
  wire       [7:0]    pes_11_10_io_outputB;
  wire       [19:0]   pes_11_10_io_outputC;
  wire       [7:0]    pes_11_11_io_outputA;
  wire       [7:0]    pes_11_11_io_outputB;
  wire       [19:0]   pes_11_11_io_outputC;
  wire       [7:0]    pes_11_12_io_outputA;
  wire       [7:0]    pes_11_12_io_outputB;
  wire       [19:0]   pes_11_12_io_outputC;
  wire       [7:0]    pes_11_13_io_outputA;
  wire       [7:0]    pes_11_13_io_outputB;
  wire       [19:0]   pes_11_13_io_outputC;
  wire       [7:0]    pes_11_14_io_outputA;
  wire       [7:0]    pes_11_14_io_outputB;
  wire       [19:0]   pes_11_14_io_outputC;
  wire       [7:0]    pes_11_15_io_outputB;
  wire       [19:0]   pes_11_15_io_outputC;
  wire       [7:0]    pes_12_0_io_outputA;
  wire       [7:0]    pes_12_0_io_outputB;
  wire       [19:0]   pes_12_0_io_outputC;
  wire       [7:0]    pes_12_1_io_outputA;
  wire       [7:0]    pes_12_1_io_outputB;
  wire       [19:0]   pes_12_1_io_outputC;
  wire       [7:0]    pes_12_2_io_outputA;
  wire       [7:0]    pes_12_2_io_outputB;
  wire       [19:0]   pes_12_2_io_outputC;
  wire       [7:0]    pes_12_3_io_outputA;
  wire       [7:0]    pes_12_3_io_outputB;
  wire       [19:0]   pes_12_3_io_outputC;
  wire       [7:0]    pes_12_4_io_outputA;
  wire       [7:0]    pes_12_4_io_outputB;
  wire       [19:0]   pes_12_4_io_outputC;
  wire       [7:0]    pes_12_5_io_outputA;
  wire       [7:0]    pes_12_5_io_outputB;
  wire       [19:0]   pes_12_5_io_outputC;
  wire       [7:0]    pes_12_6_io_outputA;
  wire       [7:0]    pes_12_6_io_outputB;
  wire       [19:0]   pes_12_6_io_outputC;
  wire       [7:0]    pes_12_7_io_outputA;
  wire       [7:0]    pes_12_7_io_outputB;
  wire       [19:0]   pes_12_7_io_outputC;
  wire       [7:0]    pes_12_8_io_outputA;
  wire       [7:0]    pes_12_8_io_outputB;
  wire       [19:0]   pes_12_8_io_outputC;
  wire       [7:0]    pes_12_9_io_outputA;
  wire       [7:0]    pes_12_9_io_outputB;
  wire       [19:0]   pes_12_9_io_outputC;
  wire       [7:0]    pes_12_10_io_outputA;
  wire       [7:0]    pes_12_10_io_outputB;
  wire       [19:0]   pes_12_10_io_outputC;
  wire       [7:0]    pes_12_11_io_outputA;
  wire       [7:0]    pes_12_11_io_outputB;
  wire       [19:0]   pes_12_11_io_outputC;
  wire       [7:0]    pes_12_12_io_outputA;
  wire       [7:0]    pes_12_12_io_outputB;
  wire       [19:0]   pes_12_12_io_outputC;
  wire       [7:0]    pes_12_13_io_outputA;
  wire       [7:0]    pes_12_13_io_outputB;
  wire       [19:0]   pes_12_13_io_outputC;
  wire       [7:0]    pes_12_14_io_outputA;
  wire       [7:0]    pes_12_14_io_outputB;
  wire       [19:0]   pes_12_14_io_outputC;
  wire       [7:0]    pes_12_15_io_outputB;
  wire       [19:0]   pes_12_15_io_outputC;
  wire       [7:0]    pes_13_0_io_outputA;
  wire       [7:0]    pes_13_0_io_outputB;
  wire       [19:0]   pes_13_0_io_outputC;
  wire       [7:0]    pes_13_1_io_outputA;
  wire       [7:0]    pes_13_1_io_outputB;
  wire       [19:0]   pes_13_1_io_outputC;
  wire       [7:0]    pes_13_2_io_outputA;
  wire       [7:0]    pes_13_2_io_outputB;
  wire       [19:0]   pes_13_2_io_outputC;
  wire       [7:0]    pes_13_3_io_outputA;
  wire       [7:0]    pes_13_3_io_outputB;
  wire       [19:0]   pes_13_3_io_outputC;
  wire       [7:0]    pes_13_4_io_outputA;
  wire       [7:0]    pes_13_4_io_outputB;
  wire       [19:0]   pes_13_4_io_outputC;
  wire       [7:0]    pes_13_5_io_outputA;
  wire       [7:0]    pes_13_5_io_outputB;
  wire       [19:0]   pes_13_5_io_outputC;
  wire       [7:0]    pes_13_6_io_outputA;
  wire       [7:0]    pes_13_6_io_outputB;
  wire       [19:0]   pes_13_6_io_outputC;
  wire       [7:0]    pes_13_7_io_outputA;
  wire       [7:0]    pes_13_7_io_outputB;
  wire       [19:0]   pes_13_7_io_outputC;
  wire       [7:0]    pes_13_8_io_outputA;
  wire       [7:0]    pes_13_8_io_outputB;
  wire       [19:0]   pes_13_8_io_outputC;
  wire       [7:0]    pes_13_9_io_outputA;
  wire       [7:0]    pes_13_9_io_outputB;
  wire       [19:0]   pes_13_9_io_outputC;
  wire       [7:0]    pes_13_10_io_outputA;
  wire       [7:0]    pes_13_10_io_outputB;
  wire       [19:0]   pes_13_10_io_outputC;
  wire       [7:0]    pes_13_11_io_outputA;
  wire       [7:0]    pes_13_11_io_outputB;
  wire       [19:0]   pes_13_11_io_outputC;
  wire       [7:0]    pes_13_12_io_outputA;
  wire       [7:0]    pes_13_12_io_outputB;
  wire       [19:0]   pes_13_12_io_outputC;
  wire       [7:0]    pes_13_13_io_outputA;
  wire       [7:0]    pes_13_13_io_outputB;
  wire       [19:0]   pes_13_13_io_outputC;
  wire       [7:0]    pes_13_14_io_outputA;
  wire       [7:0]    pes_13_14_io_outputB;
  wire       [19:0]   pes_13_14_io_outputC;
  wire       [7:0]    pes_13_15_io_outputB;
  wire       [19:0]   pes_13_15_io_outputC;
  wire       [7:0]    pes_14_0_io_outputA;
  wire       [7:0]    pes_14_0_io_outputB;
  wire       [19:0]   pes_14_0_io_outputC;
  wire       [7:0]    pes_14_1_io_outputA;
  wire       [7:0]    pes_14_1_io_outputB;
  wire       [19:0]   pes_14_1_io_outputC;
  wire       [7:0]    pes_14_2_io_outputA;
  wire       [7:0]    pes_14_2_io_outputB;
  wire       [19:0]   pes_14_2_io_outputC;
  wire       [7:0]    pes_14_3_io_outputA;
  wire       [7:0]    pes_14_3_io_outputB;
  wire       [19:0]   pes_14_3_io_outputC;
  wire       [7:0]    pes_14_4_io_outputA;
  wire       [7:0]    pes_14_4_io_outputB;
  wire       [19:0]   pes_14_4_io_outputC;
  wire       [7:0]    pes_14_5_io_outputA;
  wire       [7:0]    pes_14_5_io_outputB;
  wire       [19:0]   pes_14_5_io_outputC;
  wire       [7:0]    pes_14_6_io_outputA;
  wire       [7:0]    pes_14_6_io_outputB;
  wire       [19:0]   pes_14_6_io_outputC;
  wire       [7:0]    pes_14_7_io_outputA;
  wire       [7:0]    pes_14_7_io_outputB;
  wire       [19:0]   pes_14_7_io_outputC;
  wire       [7:0]    pes_14_8_io_outputA;
  wire       [7:0]    pes_14_8_io_outputB;
  wire       [19:0]   pes_14_8_io_outputC;
  wire       [7:0]    pes_14_9_io_outputA;
  wire       [7:0]    pes_14_9_io_outputB;
  wire       [19:0]   pes_14_9_io_outputC;
  wire       [7:0]    pes_14_10_io_outputA;
  wire       [7:0]    pes_14_10_io_outputB;
  wire       [19:0]   pes_14_10_io_outputC;
  wire       [7:0]    pes_14_11_io_outputA;
  wire       [7:0]    pes_14_11_io_outputB;
  wire       [19:0]   pes_14_11_io_outputC;
  wire       [7:0]    pes_14_12_io_outputA;
  wire       [7:0]    pes_14_12_io_outputB;
  wire       [19:0]   pes_14_12_io_outputC;
  wire       [7:0]    pes_14_13_io_outputA;
  wire       [7:0]    pes_14_13_io_outputB;
  wire       [19:0]   pes_14_13_io_outputC;
  wire       [7:0]    pes_14_14_io_outputA;
  wire       [7:0]    pes_14_14_io_outputB;
  wire       [19:0]   pes_14_14_io_outputC;
  wire       [7:0]    pes_14_15_io_outputB;
  wire       [19:0]   pes_14_15_io_outputC;
  wire       [7:0]    pes_15_0_io_outputA;
  wire       [19:0]   pes_15_0_io_outputC;
  wire       [7:0]    pes_15_1_io_outputA;
  wire       [19:0]   pes_15_1_io_outputC;
  wire       [7:0]    pes_15_2_io_outputA;
  wire       [19:0]   pes_15_2_io_outputC;
  wire       [7:0]    pes_15_3_io_outputA;
  wire       [19:0]   pes_15_3_io_outputC;
  wire       [7:0]    pes_15_4_io_outputA;
  wire       [19:0]   pes_15_4_io_outputC;
  wire       [7:0]    pes_15_5_io_outputA;
  wire       [19:0]   pes_15_5_io_outputC;
  wire       [7:0]    pes_15_6_io_outputA;
  wire       [19:0]   pes_15_6_io_outputC;
  wire       [7:0]    pes_15_7_io_outputA;
  wire       [19:0]   pes_15_7_io_outputC;
  wire       [7:0]    pes_15_8_io_outputA;
  wire       [19:0]   pes_15_8_io_outputC;
  wire       [7:0]    pes_15_9_io_outputA;
  wire       [19:0]   pes_15_9_io_outputC;
  wire       [7:0]    pes_15_10_io_outputA;
  wire       [19:0]   pes_15_10_io_outputC;
  wire       [7:0]    pes_15_11_io_outputA;
  wire       [19:0]   pes_15_11_io_outputC;
  wire       [7:0]    pes_15_12_io_outputA;
  wire       [19:0]   pes_15_12_io_outputC;
  wire       [7:0]    pes_15_13_io_outputA;
  wire       [19:0]   pes_15_13_io_outputC;
  wire       [7:0]    pes_15_14_io_outputA;
  wire       [19:0]   pes_15_14_io_outputC;
  wire       [19:0]   pes_15_15_io_outputC;
  wire       [7:0]    skewBuffer_io_output_0;
  wire       [7:0]    skewBuffer_io_output_1;
  wire       [7:0]    skewBuffer_io_output_2;
  wire       [7:0]    skewBuffer_io_output_3;
  wire       [7:0]    skewBuffer_io_output_4;
  wire       [7:0]    skewBuffer_io_output_5;
  wire       [7:0]    skewBuffer_io_output_6;
  wire       [7:0]    skewBuffer_io_output_7;
  wire       [7:0]    skewBuffer_io_output_8;
  wire       [7:0]    skewBuffer_io_output_9;
  wire       [7:0]    skewBuffer_io_output_10;
  wire       [7:0]    skewBuffer_io_output_11;
  wire       [7:0]    skewBuffer_io_output_12;
  wire       [7:0]    skewBuffer_io_output_13;
  wire       [7:0]    skewBuffer_io_output_14;
  wire       [7:0]    skewBuffer_io_output_15;
  wire       [19:0]   skewBuffer_1_io_output_0;
  wire       [19:0]   skewBuffer_1_io_output_1;
  wire       [19:0]   skewBuffer_1_io_output_2;
  wire       [19:0]   skewBuffer_1_io_output_3;
  wire       [19:0]   skewBuffer_1_io_output_4;
  wire       [19:0]   skewBuffer_1_io_output_5;
  wire       [19:0]   skewBuffer_1_io_output_6;
  wire       [19:0]   skewBuffer_1_io_output_7;
  wire       [19:0]   skewBuffer_1_io_output_8;
  wire       [19:0]   skewBuffer_1_io_output_9;
  wire       [19:0]   skewBuffer_1_io_output_10;
  wire       [19:0]   skewBuffer_1_io_output_11;
  wire       [19:0]   skewBuffer_1_io_output_12;
  wire       [19:0]   skewBuffer_1_io_output_13;
  wire       [19:0]   skewBuffer_1_io_output_14;
  wire       [19:0]   skewBuffer_1_io_output_15;
  reg        [7:0]    io_inputB_0_regNext;
  reg        [7:0]    io_inputB_1_regNext;
  reg        [7:0]    io_inputB_2_regNext;
  reg        [7:0]    io_inputB_3_regNext;
  reg        [7:0]    io_inputB_4_regNext;
  reg        [7:0]    io_inputB_5_regNext;
  reg        [7:0]    io_inputB_6_regNext;
  reg        [7:0]    io_inputB_7_regNext;
  reg        [7:0]    io_inputB_8_regNext;
  reg        [7:0]    io_inputB_9_regNext;
  reg        [7:0]    io_inputB_10_regNext;
  reg        [7:0]    io_inputB_11_regNext;
  reg        [7:0]    io_inputB_12_regNext;
  reg        [7:0]    io_inputB_13_regNext;
  reg        [7:0]    io_inputB_14_regNext;
  reg        [7:0]    io_inputB_15_regNext;
//#endregion

//#region Processing Elements
  ProcessingElement pes_0_0 (
    .io_inputA              (skewBuffer_io_output_0[7:0]), //i
    .io_inputB              (io_inputB_0_regNext[7:0]   ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_0_0 ), //i
    .io_outputA             (pes_0_0_io_outputA[7:0]    ), //o
    .io_outputB             (pes_0_0_io_outputB[7:0]    ), //o
    .io_outputC             (pes_0_0_io_outputC[15:0]   ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement pes_0_1 (
    .io_inputA              (pes_0_0_io_outputA[7:0]   ), //i
    .io_inputB              (io_inputB_1_regNext[7:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_0_1), //i
    .io_outputA             (pes_0_1_io_outputA[7:0]   ), //o
    .io_outputB             (pes_0_1_io_outputB[7:0]   ), //o
    .io_outputC             (pes_0_1_io_outputC[15:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement pes_0_2 (
    .io_inputA              (pes_0_1_io_outputA[7:0]   ), //i
    .io_inputB              (io_inputB_2_regNext[7:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_0_2), //i
    .io_outputA             (pes_0_2_io_outputA[7:0]   ), //o
    .io_outputB             (pes_0_2_io_outputB[7:0]   ), //o
    .io_outputC             (pes_0_2_io_outputC[15:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement pes_0_3 (
    .io_inputA              (pes_0_2_io_outputA[7:0]   ), //i
    .io_inputB              (io_inputB_3_regNext[7:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_0_3), //i
    .io_outputA             (pes_0_3_io_outputA[7:0]   ), //o
    .io_outputB             (pes_0_3_io_outputB[7:0]   ), //o
    .io_outputC             (pes_0_3_io_outputC[15:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement pes_0_4 (
    .io_inputA              (pes_0_3_io_outputA[7:0]   ), //i
    .io_inputB              (io_inputB_4_regNext[7:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_0_4), //i
    .io_outputA             (pes_0_4_io_outputA[7:0]   ), //o
    .io_outputB             (pes_0_4_io_outputB[7:0]   ), //o
    .io_outputC             (pes_0_4_io_outputC[15:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement pes_0_5 (
    .io_inputA              (pes_0_4_io_outputA[7:0]   ), //i
    .io_inputB              (io_inputB_5_regNext[7:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_0_5), //i
    .io_outputA             (pes_0_5_io_outputA[7:0]   ), //o
    .io_outputB             (pes_0_5_io_outputB[7:0]   ), //o
    .io_outputC             (pes_0_5_io_outputC[15:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement pes_0_6 (
    .io_inputA              (pes_0_5_io_outputA[7:0]   ), //i
    .io_inputB              (io_inputB_6_regNext[7:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_0_6), //i
    .io_outputA             (pes_0_6_io_outputA[7:0]   ), //o
    .io_outputB             (pes_0_6_io_outputB[7:0]   ), //o
    .io_outputC             (pes_0_6_io_outputC[15:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement pes_0_7 (
    .io_inputA              (pes_0_6_io_outputA[7:0]   ), //i
    .io_inputB              (io_inputB_7_regNext[7:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_0_7), //i
    .io_outputA             (pes_0_7_io_outputA[7:0]   ), //o
    .io_outputB             (pes_0_7_io_outputB[7:0]   ), //o
    .io_outputC             (pes_0_7_io_outputC[15:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement pes_0_8 (
    .io_inputA              (pes_0_7_io_outputA[7:0]   ), //i
    .io_inputB              (io_inputB_8_regNext[7:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_0_8), //i
    .io_outputA             (pes_0_8_io_outputA[7:0]   ), //o
    .io_outputB             (pes_0_8_io_outputB[7:0]   ), //o
    .io_outputC             (pes_0_8_io_outputC[15:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement pes_0_9 (
    .io_inputA              (pes_0_8_io_outputA[7:0]   ), //i
    .io_inputB              (io_inputB_9_regNext[7:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_0_9), //i
    .io_outputA             (pes_0_9_io_outputA[7:0]   ), //o
    .io_outputB             (pes_0_9_io_outputB[7:0]   ), //o
    .io_outputC             (pes_0_9_io_outputC[15:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement pes_0_10 (
    .io_inputA              (pes_0_9_io_outputA[7:0]    ), //i
    .io_inputB              (io_inputB_10_regNext[7:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_0_10), //i
    .io_outputA             (pes_0_10_io_outputA[7:0]   ), //o
    .io_outputB             (pes_0_10_io_outputB[7:0]   ), //o
    .io_outputC             (pes_0_10_io_outputC[15:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement pes_0_11 (
    .io_inputA              (pes_0_10_io_outputA[7:0]   ), //i
    .io_inputB              (io_inputB_11_regNext[7:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_0_11), //i
    .io_outputA             (pes_0_11_io_outputA[7:0]   ), //o
    .io_outputB             (pes_0_11_io_outputB[7:0]   ), //o
    .io_outputC             (pes_0_11_io_outputC[15:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement pes_0_12 (
    .io_inputA              (pes_0_11_io_outputA[7:0]   ), //i
    .io_inputB              (io_inputB_12_regNext[7:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_0_12), //i
    .io_outputA             (pes_0_12_io_outputA[7:0]   ), //o
    .io_outputB             (pes_0_12_io_outputB[7:0]   ), //o
    .io_outputC             (pes_0_12_io_outputC[15:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement pes_0_13 (
    .io_inputA              (pes_0_12_io_outputA[7:0]   ), //i
    .io_inputB              (io_inputB_13_regNext[7:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_0_13), //i
    .io_outputA             (pes_0_13_io_outputA[7:0]   ), //o
    .io_outputB             (pes_0_13_io_outputB[7:0]   ), //o
    .io_outputC             (pes_0_13_io_outputC[15:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement pes_0_14 (
    .io_inputA              (pes_0_13_io_outputA[7:0]   ), //i
    .io_inputB              (io_inputB_14_regNext[7:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_0_14), //i
    .io_outputA             (pes_0_14_io_outputA[7:0]   ), //o
    .io_outputB             (pes_0_14_io_outputB[7:0]   ), //o
    .io_outputC             (pes_0_14_io_outputC[15:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_15 pes_0_15 (
    .io_inputA              (pes_0_14_io_outputA[7:0]   ), //i
    .io_inputB              (io_inputB_15_regNext[7:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_0_15), //i
    .io_outputB             (pes_0_15_io_outputB[7:0]   ), //o
    .io_outputC             (pes_0_15_io_outputC[15:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_16 pes_1_0 (
    .io_inputA              (skewBuffer_io_output_1[7:0]), //i
    .io_inputB              (pes_0_0_io_outputB[7:0]    ), //i
    .io_inputC              (pes_0_0_io_outputC[15:0]   ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_1_0 ), //i
    .io_outputA             (pes_1_0_io_outputA[7:0]    ), //o
    .io_outputB             (pes_1_0_io_outputB[7:0]    ), //o
    .io_outputC             (pes_1_0_io_outputC[16:0]   ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_16 pes_1_1 (
    .io_inputA              (pes_1_0_io_outputA[7:0]   ), //i
    .io_inputB              (pes_0_1_io_outputB[7:0]   ), //i
    .io_inputC              (pes_0_1_io_outputC[15:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_1_1), //i
    .io_outputA             (pes_1_1_io_outputA[7:0]   ), //o
    .io_outputB             (pes_1_1_io_outputB[7:0]   ), //o
    .io_outputC             (pes_1_1_io_outputC[16:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement_16 pes_1_2 (
    .io_inputA              (pes_1_1_io_outputA[7:0]   ), //i
    .io_inputB              (pes_0_2_io_outputB[7:0]   ), //i
    .io_inputC              (pes_0_2_io_outputC[15:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_1_2), //i
    .io_outputA             (pes_1_2_io_outputA[7:0]   ), //o
    .io_outputB             (pes_1_2_io_outputB[7:0]   ), //o
    .io_outputC             (pes_1_2_io_outputC[16:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement_16 pes_1_3 (
    .io_inputA              (pes_1_2_io_outputA[7:0]   ), //i
    .io_inputB              (pes_0_3_io_outputB[7:0]   ), //i
    .io_inputC              (pes_0_3_io_outputC[15:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_1_3), //i
    .io_outputA             (pes_1_3_io_outputA[7:0]   ), //o
    .io_outputB             (pes_1_3_io_outputB[7:0]   ), //o
    .io_outputC             (pes_1_3_io_outputC[16:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement_16 pes_1_4 (
    .io_inputA              (pes_1_3_io_outputA[7:0]   ), //i
    .io_inputB              (pes_0_4_io_outputB[7:0]   ), //i
    .io_inputC              (pes_0_4_io_outputC[15:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_1_4), //i
    .io_outputA             (pes_1_4_io_outputA[7:0]   ), //o
    .io_outputB             (pes_1_4_io_outputB[7:0]   ), //o
    .io_outputC             (pes_1_4_io_outputC[16:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement_16 pes_1_5 (
    .io_inputA              (pes_1_4_io_outputA[7:0]   ), //i
    .io_inputB              (pes_0_5_io_outputB[7:0]   ), //i
    .io_inputC              (pes_0_5_io_outputC[15:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_1_5), //i
    .io_outputA             (pes_1_5_io_outputA[7:0]   ), //o
    .io_outputB             (pes_1_5_io_outputB[7:0]   ), //o
    .io_outputC             (pes_1_5_io_outputC[16:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement_16 pes_1_6 (
    .io_inputA              (pes_1_5_io_outputA[7:0]   ), //i
    .io_inputB              (pes_0_6_io_outputB[7:0]   ), //i
    .io_inputC              (pes_0_6_io_outputC[15:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_1_6), //i
    .io_outputA             (pes_1_6_io_outputA[7:0]   ), //o
    .io_outputB             (pes_1_6_io_outputB[7:0]   ), //o
    .io_outputC             (pes_1_6_io_outputC[16:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement_16 pes_1_7 (
    .io_inputA              (pes_1_6_io_outputA[7:0]   ), //i
    .io_inputB              (pes_0_7_io_outputB[7:0]   ), //i
    .io_inputC              (pes_0_7_io_outputC[15:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_1_7), //i
    .io_outputA             (pes_1_7_io_outputA[7:0]   ), //o
    .io_outputB             (pes_1_7_io_outputB[7:0]   ), //o
    .io_outputC             (pes_1_7_io_outputC[16:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement_16 pes_1_8 (
    .io_inputA              (pes_1_7_io_outputA[7:0]   ), //i
    .io_inputB              (pes_0_8_io_outputB[7:0]   ), //i
    .io_inputC              (pes_0_8_io_outputC[15:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_1_8), //i
    .io_outputA             (pes_1_8_io_outputA[7:0]   ), //o
    .io_outputB             (pes_1_8_io_outputB[7:0]   ), //o
    .io_outputC             (pes_1_8_io_outputC[16:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement_16 pes_1_9 (
    .io_inputA              (pes_1_8_io_outputA[7:0]   ), //i
    .io_inputB              (pes_0_9_io_outputB[7:0]   ), //i
    .io_inputC              (pes_0_9_io_outputC[15:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_1_9), //i
    .io_outputA             (pes_1_9_io_outputA[7:0]   ), //o
    .io_outputB             (pes_1_9_io_outputB[7:0]   ), //o
    .io_outputC             (pes_1_9_io_outputC[16:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement_16 pes_1_10 (
    .io_inputA              (pes_1_9_io_outputA[7:0]    ), //i
    .io_inputB              (pes_0_10_io_outputB[7:0]   ), //i
    .io_inputC              (pes_0_10_io_outputC[15:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_1_10), //i
    .io_outputA             (pes_1_10_io_outputA[7:0]   ), //o
    .io_outputB             (pes_1_10_io_outputB[7:0]   ), //o
    .io_outputC             (pes_1_10_io_outputC[16:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_16 pes_1_11 (
    .io_inputA              (pes_1_10_io_outputA[7:0]   ), //i
    .io_inputB              (pes_0_11_io_outputB[7:0]   ), //i
    .io_inputC              (pes_0_11_io_outputC[15:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_1_11), //i
    .io_outputA             (pes_1_11_io_outputA[7:0]   ), //o
    .io_outputB             (pes_1_11_io_outputB[7:0]   ), //o
    .io_outputC             (pes_1_11_io_outputC[16:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_16 pes_1_12 (
    .io_inputA              (pes_1_11_io_outputA[7:0]   ), //i
    .io_inputB              (pes_0_12_io_outputB[7:0]   ), //i
    .io_inputC              (pes_0_12_io_outputC[15:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_1_12), //i
    .io_outputA             (pes_1_12_io_outputA[7:0]   ), //o
    .io_outputB             (pes_1_12_io_outputB[7:0]   ), //o
    .io_outputC             (pes_1_12_io_outputC[16:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_16 pes_1_13 (
    .io_inputA              (pes_1_12_io_outputA[7:0]   ), //i
    .io_inputB              (pes_0_13_io_outputB[7:0]   ), //i
    .io_inputC              (pes_0_13_io_outputC[15:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_1_13), //i
    .io_outputA             (pes_1_13_io_outputA[7:0]   ), //o
    .io_outputB             (pes_1_13_io_outputB[7:0]   ), //o
    .io_outputC             (pes_1_13_io_outputC[16:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_16 pes_1_14 (
    .io_inputA              (pes_1_13_io_outputA[7:0]   ), //i
    .io_inputB              (pes_0_14_io_outputB[7:0]   ), //i
    .io_inputC              (pes_0_14_io_outputC[15:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_1_14), //i
    .io_outputA             (pes_1_14_io_outputA[7:0]   ), //o
    .io_outputB             (pes_1_14_io_outputB[7:0]   ), //o
    .io_outputC             (pes_1_14_io_outputC[16:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_31 pes_1_15 (
    .io_inputA              (pes_1_14_io_outputA[7:0]   ), //i
    .io_inputB              (pes_0_15_io_outputB[7:0]   ), //i
    .io_inputC              (pes_0_15_io_outputC[15:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_1_15), //i
    .io_outputB             (pes_1_15_io_outputB[7:0]   ), //o
    .io_outputC             (pes_1_15_io_outputC[16:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_32 pes_2_0 (
    .io_inputA              (skewBuffer_io_output_2[7:0]), //i
    .io_inputB              (pes_1_0_io_outputB[7:0]    ), //i
    .io_inputC              (pes_1_0_io_outputC[16:0]   ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_2_0 ), //i
    .io_outputA             (pes_2_0_io_outputA[7:0]    ), //o
    .io_outputB             (pes_2_0_io_outputB[7:0]    ), //o
    .io_outputC             (pes_2_0_io_outputC[17:0]   ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_32 pes_2_1 (
    .io_inputA              (pes_2_0_io_outputA[7:0]   ), //i
    .io_inputB              (pes_1_1_io_outputB[7:0]   ), //i
    .io_inputC              (pes_1_1_io_outputC[16:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_2_1), //i
    .io_outputA             (pes_2_1_io_outputA[7:0]   ), //o
    .io_outputB             (pes_2_1_io_outputB[7:0]   ), //o
    .io_outputC             (pes_2_1_io_outputC[17:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement_32 pes_2_2 (
    .io_inputA              (pes_2_1_io_outputA[7:0]   ), //i
    .io_inputB              (pes_1_2_io_outputB[7:0]   ), //i
    .io_inputC              (pes_1_2_io_outputC[16:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_2_2), //i
    .io_outputA             (pes_2_2_io_outputA[7:0]   ), //o
    .io_outputB             (pes_2_2_io_outputB[7:0]   ), //o
    .io_outputC             (pes_2_2_io_outputC[17:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement_32 pes_2_3 (
    .io_inputA              (pes_2_2_io_outputA[7:0]   ), //i
    .io_inputB              (pes_1_3_io_outputB[7:0]   ), //i
    .io_inputC              (pes_1_3_io_outputC[16:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_2_3), //i
    .io_outputA             (pes_2_3_io_outputA[7:0]   ), //o
    .io_outputB             (pes_2_3_io_outputB[7:0]   ), //o
    .io_outputC             (pes_2_3_io_outputC[17:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement_32 pes_2_4 (
    .io_inputA              (pes_2_3_io_outputA[7:0]   ), //i
    .io_inputB              (pes_1_4_io_outputB[7:0]   ), //i
    .io_inputC              (pes_1_4_io_outputC[16:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_2_4), //i
    .io_outputA             (pes_2_4_io_outputA[7:0]   ), //o
    .io_outputB             (pes_2_4_io_outputB[7:0]   ), //o
    .io_outputC             (pes_2_4_io_outputC[17:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement_32 pes_2_5 (
    .io_inputA              (pes_2_4_io_outputA[7:0]   ), //i
    .io_inputB              (pes_1_5_io_outputB[7:0]   ), //i
    .io_inputC              (pes_1_5_io_outputC[16:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_2_5), //i
    .io_outputA             (pes_2_5_io_outputA[7:0]   ), //o
    .io_outputB             (pes_2_5_io_outputB[7:0]   ), //o
    .io_outputC             (pes_2_5_io_outputC[17:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement_32 pes_2_6 (
    .io_inputA              (pes_2_5_io_outputA[7:0]   ), //i
    .io_inputB              (pes_1_6_io_outputB[7:0]   ), //i
    .io_inputC              (pes_1_6_io_outputC[16:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_2_6), //i
    .io_outputA             (pes_2_6_io_outputA[7:0]   ), //o
    .io_outputB             (pes_2_6_io_outputB[7:0]   ), //o
    .io_outputC             (pes_2_6_io_outputC[17:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement_32 pes_2_7 (
    .io_inputA              (pes_2_6_io_outputA[7:0]   ), //i
    .io_inputB              (pes_1_7_io_outputB[7:0]   ), //i
    .io_inputC              (pes_1_7_io_outputC[16:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_2_7), //i
    .io_outputA             (pes_2_7_io_outputA[7:0]   ), //o
    .io_outputB             (pes_2_7_io_outputB[7:0]   ), //o
    .io_outputC             (pes_2_7_io_outputC[17:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement_32 pes_2_8 (
    .io_inputA              (pes_2_7_io_outputA[7:0]   ), //i
    .io_inputB              (pes_1_8_io_outputB[7:0]   ), //i
    .io_inputC              (pes_1_8_io_outputC[16:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_2_8), //i
    .io_outputA             (pes_2_8_io_outputA[7:0]   ), //o
    .io_outputB             (pes_2_8_io_outputB[7:0]   ), //o
    .io_outputC             (pes_2_8_io_outputC[17:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement_32 pes_2_9 (
    .io_inputA              (pes_2_8_io_outputA[7:0]   ), //i
    .io_inputB              (pes_1_9_io_outputB[7:0]   ), //i
    .io_inputC              (pes_1_9_io_outputC[16:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_2_9), //i
    .io_outputA             (pes_2_9_io_outputA[7:0]   ), //o
    .io_outputB             (pes_2_9_io_outputB[7:0]   ), //o
    .io_outputC             (pes_2_9_io_outputC[17:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement_32 pes_2_10 (
    .io_inputA              (pes_2_9_io_outputA[7:0]    ), //i
    .io_inputB              (pes_1_10_io_outputB[7:0]   ), //i
    .io_inputC              (pes_1_10_io_outputC[16:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_2_10), //i
    .io_outputA             (pes_2_10_io_outputA[7:0]   ), //o
    .io_outputB             (pes_2_10_io_outputB[7:0]   ), //o
    .io_outputC             (pes_2_10_io_outputC[17:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_32 pes_2_11 (
    .io_inputA              (pes_2_10_io_outputA[7:0]   ), //i
    .io_inputB              (pes_1_11_io_outputB[7:0]   ), //i
    .io_inputC              (pes_1_11_io_outputC[16:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_2_11), //i
    .io_outputA             (pes_2_11_io_outputA[7:0]   ), //o
    .io_outputB             (pes_2_11_io_outputB[7:0]   ), //o
    .io_outputC             (pes_2_11_io_outputC[17:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_32 pes_2_12 (
    .io_inputA              (pes_2_11_io_outputA[7:0]   ), //i
    .io_inputB              (pes_1_12_io_outputB[7:0]   ), //i
    .io_inputC              (pes_1_12_io_outputC[16:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_2_12), //i
    .io_outputA             (pes_2_12_io_outputA[7:0]   ), //o
    .io_outputB             (pes_2_12_io_outputB[7:0]   ), //o
    .io_outputC             (pes_2_12_io_outputC[17:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_32 pes_2_13 (
    .io_inputA              (pes_2_12_io_outputA[7:0]   ), //i
    .io_inputB              (pes_1_13_io_outputB[7:0]   ), //i
    .io_inputC              (pes_1_13_io_outputC[16:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_2_13), //i
    .io_outputA             (pes_2_13_io_outputA[7:0]   ), //o
    .io_outputB             (pes_2_13_io_outputB[7:0]   ), //o
    .io_outputC             (pes_2_13_io_outputC[17:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_32 pes_2_14 (
    .io_inputA              (pes_2_13_io_outputA[7:0]   ), //i
    .io_inputB              (pes_1_14_io_outputB[7:0]   ), //i
    .io_inputC              (pes_1_14_io_outputC[16:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_2_14), //i
    .io_outputA             (pes_2_14_io_outputA[7:0]   ), //o
    .io_outputB             (pes_2_14_io_outputB[7:0]   ), //o
    .io_outputC             (pes_2_14_io_outputC[17:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_47 pes_2_15 (
    .io_inputA              (pes_2_14_io_outputA[7:0]   ), //i
    .io_inputB              (pes_1_15_io_outputB[7:0]   ), //i
    .io_inputC              (pes_1_15_io_outputC[16:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_2_15), //i
    .io_outputB             (pes_2_15_io_outputB[7:0]   ), //o
    .io_outputC             (pes_2_15_io_outputC[17:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_48 pes_3_0 (
    .io_inputA              (skewBuffer_io_output_3[7:0]), //i
    .io_inputB              (pes_2_0_io_outputB[7:0]    ), //i
    .io_inputC              (pes_2_0_io_outputC[17:0]   ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_3_0 ), //i
    .io_outputA             (pes_3_0_io_outputA[7:0]    ), //o
    .io_outputB             (pes_3_0_io_outputB[7:0]    ), //o
    .io_outputC             (pes_3_0_io_outputC[17:0]   ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_48 pes_3_1 (
    .io_inputA              (pes_3_0_io_outputA[7:0]   ), //i
    .io_inputB              (pes_2_1_io_outputB[7:0]   ), //i
    .io_inputC              (pes_2_1_io_outputC[17:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_3_1), //i
    .io_outputA             (pes_3_1_io_outputA[7:0]   ), //o
    .io_outputB             (pes_3_1_io_outputB[7:0]   ), //o
    .io_outputC             (pes_3_1_io_outputC[17:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement_48 pes_3_2 (
    .io_inputA              (pes_3_1_io_outputA[7:0]   ), //i
    .io_inputB              (pes_2_2_io_outputB[7:0]   ), //i
    .io_inputC              (pes_2_2_io_outputC[17:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_3_2), //i
    .io_outputA             (pes_3_2_io_outputA[7:0]   ), //o
    .io_outputB             (pes_3_2_io_outputB[7:0]   ), //o
    .io_outputC             (pes_3_2_io_outputC[17:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement_48 pes_3_3 (
    .io_inputA              (pes_3_2_io_outputA[7:0]   ), //i
    .io_inputB              (pes_2_3_io_outputB[7:0]   ), //i
    .io_inputC              (pes_2_3_io_outputC[17:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_3_3), //i
    .io_outputA             (pes_3_3_io_outputA[7:0]   ), //o
    .io_outputB             (pes_3_3_io_outputB[7:0]   ), //o
    .io_outputC             (pes_3_3_io_outputC[17:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement_48 pes_3_4 (
    .io_inputA              (pes_3_3_io_outputA[7:0]   ), //i
    .io_inputB              (pes_2_4_io_outputB[7:0]   ), //i
    .io_inputC              (pes_2_4_io_outputC[17:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_3_4), //i
    .io_outputA             (pes_3_4_io_outputA[7:0]   ), //o
    .io_outputB             (pes_3_4_io_outputB[7:0]   ), //o
    .io_outputC             (pes_3_4_io_outputC[17:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement_48 pes_3_5 (
    .io_inputA              (pes_3_4_io_outputA[7:0]   ), //i
    .io_inputB              (pes_2_5_io_outputB[7:0]   ), //i
    .io_inputC              (pes_2_5_io_outputC[17:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_3_5), //i
    .io_outputA             (pes_3_5_io_outputA[7:0]   ), //o
    .io_outputB             (pes_3_5_io_outputB[7:0]   ), //o
    .io_outputC             (pes_3_5_io_outputC[17:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement_48 pes_3_6 (
    .io_inputA              (pes_3_5_io_outputA[7:0]   ), //i
    .io_inputB              (pes_2_6_io_outputB[7:0]   ), //i
    .io_inputC              (pes_2_6_io_outputC[17:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_3_6), //i
    .io_outputA             (pes_3_6_io_outputA[7:0]   ), //o
    .io_outputB             (pes_3_6_io_outputB[7:0]   ), //o
    .io_outputC             (pes_3_6_io_outputC[17:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement_48 pes_3_7 (
    .io_inputA              (pes_3_6_io_outputA[7:0]   ), //i
    .io_inputB              (pes_2_7_io_outputB[7:0]   ), //i
    .io_inputC              (pes_2_7_io_outputC[17:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_3_7), //i
    .io_outputA             (pes_3_7_io_outputA[7:0]   ), //o
    .io_outputB             (pes_3_7_io_outputB[7:0]   ), //o
    .io_outputC             (pes_3_7_io_outputC[17:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement_48 pes_3_8 (
    .io_inputA              (pes_3_7_io_outputA[7:0]   ), //i
    .io_inputB              (pes_2_8_io_outputB[7:0]   ), //i
    .io_inputC              (pes_2_8_io_outputC[17:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_3_8), //i
    .io_outputA             (pes_3_8_io_outputA[7:0]   ), //o
    .io_outputB             (pes_3_8_io_outputB[7:0]   ), //o
    .io_outputC             (pes_3_8_io_outputC[17:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement_48 pes_3_9 (
    .io_inputA              (pes_3_8_io_outputA[7:0]   ), //i
    .io_inputB              (pes_2_9_io_outputB[7:0]   ), //i
    .io_inputC              (pes_2_9_io_outputC[17:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_3_9), //i
    .io_outputA             (pes_3_9_io_outputA[7:0]   ), //o
    .io_outputB             (pes_3_9_io_outputB[7:0]   ), //o
    .io_outputC             (pes_3_9_io_outputC[17:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement_48 pes_3_10 (
    .io_inputA              (pes_3_9_io_outputA[7:0]    ), //i
    .io_inputB              (pes_2_10_io_outputB[7:0]   ), //i
    .io_inputC              (pes_2_10_io_outputC[17:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_3_10), //i
    .io_outputA             (pes_3_10_io_outputA[7:0]   ), //o
    .io_outputB             (pes_3_10_io_outputB[7:0]   ), //o
    .io_outputC             (pes_3_10_io_outputC[17:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_48 pes_3_11 (
    .io_inputA              (pes_3_10_io_outputA[7:0]   ), //i
    .io_inputB              (pes_2_11_io_outputB[7:0]   ), //i
    .io_inputC              (pes_2_11_io_outputC[17:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_3_11), //i
    .io_outputA             (pes_3_11_io_outputA[7:0]   ), //o
    .io_outputB             (pes_3_11_io_outputB[7:0]   ), //o
    .io_outputC             (pes_3_11_io_outputC[17:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_48 pes_3_12 (
    .io_inputA              (pes_3_11_io_outputA[7:0]   ), //i
    .io_inputB              (pes_2_12_io_outputB[7:0]   ), //i
    .io_inputC              (pes_2_12_io_outputC[17:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_3_12), //i
    .io_outputA             (pes_3_12_io_outputA[7:0]   ), //o
    .io_outputB             (pes_3_12_io_outputB[7:0]   ), //o
    .io_outputC             (pes_3_12_io_outputC[17:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_48 pes_3_13 (
    .io_inputA              (pes_3_12_io_outputA[7:0]   ), //i
    .io_inputB              (pes_2_13_io_outputB[7:0]   ), //i
    .io_inputC              (pes_2_13_io_outputC[17:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_3_13), //i
    .io_outputA             (pes_3_13_io_outputA[7:0]   ), //o
    .io_outputB             (pes_3_13_io_outputB[7:0]   ), //o
    .io_outputC             (pes_3_13_io_outputC[17:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_48 pes_3_14 (
    .io_inputA              (pes_3_13_io_outputA[7:0]   ), //i
    .io_inputB              (pes_2_14_io_outputB[7:0]   ), //i
    .io_inputC              (pes_2_14_io_outputC[17:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_3_14), //i
    .io_outputA             (pes_3_14_io_outputA[7:0]   ), //o
    .io_outputB             (pes_3_14_io_outputB[7:0]   ), //o
    .io_outputC             (pes_3_14_io_outputC[17:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_63 pes_3_15 (
    .io_inputA              (pes_3_14_io_outputA[7:0]   ), //i
    .io_inputB              (pes_2_15_io_outputB[7:0]   ), //i
    .io_inputC              (pes_2_15_io_outputC[17:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_3_15), //i
    .io_outputB             (pes_3_15_io_outputB[7:0]   ), //o
    .io_outputC             (pes_3_15_io_outputC[17:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_64 pes_4_0 (
    .io_inputA              (skewBuffer_io_output_4[7:0]), //i
    .io_inputB              (pes_3_0_io_outputB[7:0]    ), //i
    .io_inputC              (pes_3_0_io_outputC[17:0]   ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_4_0 ), //i
    .io_outputA             (pes_4_0_io_outputA[7:0]    ), //o
    .io_outputB             (pes_4_0_io_outputB[7:0]    ), //o
    .io_outputC             (pes_4_0_io_outputC[18:0]   ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_64 pes_4_1 (
    .io_inputA              (pes_4_0_io_outputA[7:0]   ), //i
    .io_inputB              (pes_3_1_io_outputB[7:0]   ), //i
    .io_inputC              (pes_3_1_io_outputC[17:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_4_1), //i
    .io_outputA             (pes_4_1_io_outputA[7:0]   ), //o
    .io_outputB             (pes_4_1_io_outputB[7:0]   ), //o
    .io_outputC             (pes_4_1_io_outputC[18:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement_64 pes_4_2 (
    .io_inputA              (pes_4_1_io_outputA[7:0]   ), //i
    .io_inputB              (pes_3_2_io_outputB[7:0]   ), //i
    .io_inputC              (pes_3_2_io_outputC[17:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_4_2), //i
    .io_outputA             (pes_4_2_io_outputA[7:0]   ), //o
    .io_outputB             (pes_4_2_io_outputB[7:0]   ), //o
    .io_outputC             (pes_4_2_io_outputC[18:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement_64 pes_4_3 (
    .io_inputA              (pes_4_2_io_outputA[7:0]   ), //i
    .io_inputB              (pes_3_3_io_outputB[7:0]   ), //i
    .io_inputC              (pes_3_3_io_outputC[17:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_4_3), //i
    .io_outputA             (pes_4_3_io_outputA[7:0]   ), //o
    .io_outputB             (pes_4_3_io_outputB[7:0]   ), //o
    .io_outputC             (pes_4_3_io_outputC[18:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement_64 pes_4_4 (
    .io_inputA              (pes_4_3_io_outputA[7:0]   ), //i
    .io_inputB              (pes_3_4_io_outputB[7:0]   ), //i
    .io_inputC              (pes_3_4_io_outputC[17:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_4_4), //i
    .io_outputA             (pes_4_4_io_outputA[7:0]   ), //o
    .io_outputB             (pes_4_4_io_outputB[7:0]   ), //o
    .io_outputC             (pes_4_4_io_outputC[18:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement_64 pes_4_5 (
    .io_inputA              (pes_4_4_io_outputA[7:0]   ), //i
    .io_inputB              (pes_3_5_io_outputB[7:0]   ), //i
    .io_inputC              (pes_3_5_io_outputC[17:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_4_5), //i
    .io_outputA             (pes_4_5_io_outputA[7:0]   ), //o
    .io_outputB             (pes_4_5_io_outputB[7:0]   ), //o
    .io_outputC             (pes_4_5_io_outputC[18:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement_64 pes_4_6 (
    .io_inputA              (pes_4_5_io_outputA[7:0]   ), //i
    .io_inputB              (pes_3_6_io_outputB[7:0]   ), //i
    .io_inputC              (pes_3_6_io_outputC[17:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_4_6), //i
    .io_outputA             (pes_4_6_io_outputA[7:0]   ), //o
    .io_outputB             (pes_4_6_io_outputB[7:0]   ), //o
    .io_outputC             (pes_4_6_io_outputC[18:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement_64 pes_4_7 (
    .io_inputA              (pes_4_6_io_outputA[7:0]   ), //i
    .io_inputB              (pes_3_7_io_outputB[7:0]   ), //i
    .io_inputC              (pes_3_7_io_outputC[17:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_4_7), //i
    .io_outputA             (pes_4_7_io_outputA[7:0]   ), //o
    .io_outputB             (pes_4_7_io_outputB[7:0]   ), //o
    .io_outputC             (pes_4_7_io_outputC[18:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement_64 pes_4_8 (
    .io_inputA              (pes_4_7_io_outputA[7:0]   ), //i
    .io_inputB              (pes_3_8_io_outputB[7:0]   ), //i
    .io_inputC              (pes_3_8_io_outputC[17:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_4_8), //i
    .io_outputA             (pes_4_8_io_outputA[7:0]   ), //o
    .io_outputB             (pes_4_8_io_outputB[7:0]   ), //o
    .io_outputC             (pes_4_8_io_outputC[18:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement_64 pes_4_9 (
    .io_inputA              (pes_4_8_io_outputA[7:0]   ), //i
    .io_inputB              (pes_3_9_io_outputB[7:0]   ), //i
    .io_inputC              (pes_3_9_io_outputC[17:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_4_9), //i
    .io_outputA             (pes_4_9_io_outputA[7:0]   ), //o
    .io_outputB             (pes_4_9_io_outputB[7:0]   ), //o
    .io_outputC             (pes_4_9_io_outputC[18:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement_64 pes_4_10 (
    .io_inputA              (pes_4_9_io_outputA[7:0]    ), //i
    .io_inputB              (pes_3_10_io_outputB[7:0]   ), //i
    .io_inputC              (pes_3_10_io_outputC[17:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_4_10), //i
    .io_outputA             (pes_4_10_io_outputA[7:0]   ), //o
    .io_outputB             (pes_4_10_io_outputB[7:0]   ), //o
    .io_outputC             (pes_4_10_io_outputC[18:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_64 pes_4_11 (
    .io_inputA              (pes_4_10_io_outputA[7:0]   ), //i
    .io_inputB              (pes_3_11_io_outputB[7:0]   ), //i
    .io_inputC              (pes_3_11_io_outputC[17:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_4_11), //i
    .io_outputA             (pes_4_11_io_outputA[7:0]   ), //o
    .io_outputB             (pes_4_11_io_outputB[7:0]   ), //o
    .io_outputC             (pes_4_11_io_outputC[18:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_64 pes_4_12 (
    .io_inputA              (pes_4_11_io_outputA[7:0]   ), //i
    .io_inputB              (pes_3_12_io_outputB[7:0]   ), //i
    .io_inputC              (pes_3_12_io_outputC[17:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_4_12), //i
    .io_outputA             (pes_4_12_io_outputA[7:0]   ), //o
    .io_outputB             (pes_4_12_io_outputB[7:0]   ), //o
    .io_outputC             (pes_4_12_io_outputC[18:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_64 pes_4_13 (
    .io_inputA              (pes_4_12_io_outputA[7:0]   ), //i
    .io_inputB              (pes_3_13_io_outputB[7:0]   ), //i
    .io_inputC              (pes_3_13_io_outputC[17:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_4_13), //i
    .io_outputA             (pes_4_13_io_outputA[7:0]   ), //o
    .io_outputB             (pes_4_13_io_outputB[7:0]   ), //o
    .io_outputC             (pes_4_13_io_outputC[18:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_64 pes_4_14 (
    .io_inputA              (pes_4_13_io_outputA[7:0]   ), //i
    .io_inputB              (pes_3_14_io_outputB[7:0]   ), //i
    .io_inputC              (pes_3_14_io_outputC[17:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_4_14), //i
    .io_outputA             (pes_4_14_io_outputA[7:0]   ), //o
    .io_outputB             (pes_4_14_io_outputB[7:0]   ), //o
    .io_outputC             (pes_4_14_io_outputC[18:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_79 pes_4_15 (
    .io_inputA              (pes_4_14_io_outputA[7:0]   ), //i
    .io_inputB              (pes_3_15_io_outputB[7:0]   ), //i
    .io_inputC              (pes_3_15_io_outputC[17:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_4_15), //i
    .io_outputB             (pes_4_15_io_outputB[7:0]   ), //o
    .io_outputC             (pes_4_15_io_outputC[18:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_80 pes_5_0 (
    .io_inputA              (skewBuffer_io_output_5[7:0]), //i
    .io_inputB              (pes_4_0_io_outputB[7:0]    ), //i
    .io_inputC              (pes_4_0_io_outputC[18:0]   ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_5_0 ), //i
    .io_outputA             (pes_5_0_io_outputA[7:0]    ), //o
    .io_outputB             (pes_5_0_io_outputB[7:0]    ), //o
    .io_outputC             (pes_5_0_io_outputC[18:0]   ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_80 pes_5_1 (
    .io_inputA              (pes_5_0_io_outputA[7:0]   ), //i
    .io_inputB              (pes_4_1_io_outputB[7:0]   ), //i
    .io_inputC              (pes_4_1_io_outputC[18:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_5_1), //i
    .io_outputA             (pes_5_1_io_outputA[7:0]   ), //o
    .io_outputB             (pes_5_1_io_outputB[7:0]   ), //o
    .io_outputC             (pes_5_1_io_outputC[18:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement_80 pes_5_2 (
    .io_inputA              (pes_5_1_io_outputA[7:0]   ), //i
    .io_inputB              (pes_4_2_io_outputB[7:0]   ), //i
    .io_inputC              (pes_4_2_io_outputC[18:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_5_2), //i
    .io_outputA             (pes_5_2_io_outputA[7:0]   ), //o
    .io_outputB             (pes_5_2_io_outputB[7:0]   ), //o
    .io_outputC             (pes_5_2_io_outputC[18:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement_80 pes_5_3 (
    .io_inputA              (pes_5_2_io_outputA[7:0]   ), //i
    .io_inputB              (pes_4_3_io_outputB[7:0]   ), //i
    .io_inputC              (pes_4_3_io_outputC[18:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_5_3), //i
    .io_outputA             (pes_5_3_io_outputA[7:0]   ), //o
    .io_outputB             (pes_5_3_io_outputB[7:0]   ), //o
    .io_outputC             (pes_5_3_io_outputC[18:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement_80 pes_5_4 (
    .io_inputA              (pes_5_3_io_outputA[7:0]   ), //i
    .io_inputB              (pes_4_4_io_outputB[7:0]   ), //i
    .io_inputC              (pes_4_4_io_outputC[18:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_5_4), //i
    .io_outputA             (pes_5_4_io_outputA[7:0]   ), //o
    .io_outputB             (pes_5_4_io_outputB[7:0]   ), //o
    .io_outputC             (pes_5_4_io_outputC[18:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement_80 pes_5_5 (
    .io_inputA              (pes_5_4_io_outputA[7:0]   ), //i
    .io_inputB              (pes_4_5_io_outputB[7:0]   ), //i
    .io_inputC              (pes_4_5_io_outputC[18:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_5_5), //i
    .io_outputA             (pes_5_5_io_outputA[7:0]   ), //o
    .io_outputB             (pes_5_5_io_outputB[7:0]   ), //o
    .io_outputC             (pes_5_5_io_outputC[18:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement_80 pes_5_6 (
    .io_inputA              (pes_5_5_io_outputA[7:0]   ), //i
    .io_inputB              (pes_4_6_io_outputB[7:0]   ), //i
    .io_inputC              (pes_4_6_io_outputC[18:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_5_6), //i
    .io_outputA             (pes_5_6_io_outputA[7:0]   ), //o
    .io_outputB             (pes_5_6_io_outputB[7:0]   ), //o
    .io_outputC             (pes_5_6_io_outputC[18:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement_80 pes_5_7 (
    .io_inputA              (pes_5_6_io_outputA[7:0]   ), //i
    .io_inputB              (pes_4_7_io_outputB[7:0]   ), //i
    .io_inputC              (pes_4_7_io_outputC[18:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_5_7), //i
    .io_outputA             (pes_5_7_io_outputA[7:0]   ), //o
    .io_outputB             (pes_5_7_io_outputB[7:0]   ), //o
    .io_outputC             (pes_5_7_io_outputC[18:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement_80 pes_5_8 (
    .io_inputA              (pes_5_7_io_outputA[7:0]   ), //i
    .io_inputB              (pes_4_8_io_outputB[7:0]   ), //i
    .io_inputC              (pes_4_8_io_outputC[18:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_5_8), //i
    .io_outputA             (pes_5_8_io_outputA[7:0]   ), //o
    .io_outputB             (pes_5_8_io_outputB[7:0]   ), //o
    .io_outputC             (pes_5_8_io_outputC[18:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement_80 pes_5_9 (
    .io_inputA              (pes_5_8_io_outputA[7:0]   ), //i
    .io_inputB              (pes_4_9_io_outputB[7:0]   ), //i
    .io_inputC              (pes_4_9_io_outputC[18:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_5_9), //i
    .io_outputA             (pes_5_9_io_outputA[7:0]   ), //o
    .io_outputB             (pes_5_9_io_outputB[7:0]   ), //o
    .io_outputC             (pes_5_9_io_outputC[18:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement_80 pes_5_10 (
    .io_inputA              (pes_5_9_io_outputA[7:0]    ), //i
    .io_inputB              (pes_4_10_io_outputB[7:0]   ), //i
    .io_inputC              (pes_4_10_io_outputC[18:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_5_10), //i
    .io_outputA             (pes_5_10_io_outputA[7:0]   ), //o
    .io_outputB             (pes_5_10_io_outputB[7:0]   ), //o
    .io_outputC             (pes_5_10_io_outputC[18:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_80 pes_5_11 (
    .io_inputA              (pes_5_10_io_outputA[7:0]   ), //i
    .io_inputB              (pes_4_11_io_outputB[7:0]   ), //i
    .io_inputC              (pes_4_11_io_outputC[18:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_5_11), //i
    .io_outputA             (pes_5_11_io_outputA[7:0]   ), //o
    .io_outputB             (pes_5_11_io_outputB[7:0]   ), //o
    .io_outputC             (pes_5_11_io_outputC[18:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_80 pes_5_12 (
    .io_inputA              (pes_5_11_io_outputA[7:0]   ), //i
    .io_inputB              (pes_4_12_io_outputB[7:0]   ), //i
    .io_inputC              (pes_4_12_io_outputC[18:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_5_12), //i
    .io_outputA             (pes_5_12_io_outputA[7:0]   ), //o
    .io_outputB             (pes_5_12_io_outputB[7:0]   ), //o
    .io_outputC             (pes_5_12_io_outputC[18:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_80 pes_5_13 (
    .io_inputA              (pes_5_12_io_outputA[7:0]   ), //i
    .io_inputB              (pes_4_13_io_outputB[7:0]   ), //i
    .io_inputC              (pes_4_13_io_outputC[18:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_5_13), //i
    .io_outputA             (pes_5_13_io_outputA[7:0]   ), //o
    .io_outputB             (pes_5_13_io_outputB[7:0]   ), //o
    .io_outputC             (pes_5_13_io_outputC[18:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_80 pes_5_14 (
    .io_inputA              (pes_5_13_io_outputA[7:0]   ), //i
    .io_inputB              (pes_4_14_io_outputB[7:0]   ), //i
    .io_inputC              (pes_4_14_io_outputC[18:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_5_14), //i
    .io_outputA             (pes_5_14_io_outputA[7:0]   ), //o
    .io_outputB             (pes_5_14_io_outputB[7:0]   ), //o
    .io_outputC             (pes_5_14_io_outputC[18:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_95 pes_5_15 (
    .io_inputA              (pes_5_14_io_outputA[7:0]   ), //i
    .io_inputB              (pes_4_15_io_outputB[7:0]   ), //i
    .io_inputC              (pes_4_15_io_outputC[18:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_5_15), //i
    .io_outputB             (pes_5_15_io_outputB[7:0]   ), //o
    .io_outputC             (pes_5_15_io_outputC[18:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_80 pes_6_0 (
    .io_inputA              (skewBuffer_io_output_6[7:0]), //i
    .io_inputB              (pes_5_0_io_outputB[7:0]    ), //i
    .io_inputC              (pes_5_0_io_outputC[18:0]   ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_6_0 ), //i
    .io_outputA             (pes_6_0_io_outputA[7:0]    ), //o
    .io_outputB             (pes_6_0_io_outputB[7:0]    ), //o
    .io_outputC             (pes_6_0_io_outputC[18:0]   ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_80 pes_6_1 (
    .io_inputA              (pes_6_0_io_outputA[7:0]   ), //i
    .io_inputB              (pes_5_1_io_outputB[7:0]   ), //i
    .io_inputC              (pes_5_1_io_outputC[18:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_6_1), //i
    .io_outputA             (pes_6_1_io_outputA[7:0]   ), //o
    .io_outputB             (pes_6_1_io_outputB[7:0]   ), //o
    .io_outputC             (pes_6_1_io_outputC[18:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement_80 pes_6_2 (
    .io_inputA              (pes_6_1_io_outputA[7:0]   ), //i
    .io_inputB              (pes_5_2_io_outputB[7:0]   ), //i
    .io_inputC              (pes_5_2_io_outputC[18:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_6_2), //i
    .io_outputA             (pes_6_2_io_outputA[7:0]   ), //o
    .io_outputB             (pes_6_2_io_outputB[7:0]   ), //o
    .io_outputC             (pes_6_2_io_outputC[18:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement_80 pes_6_3 (
    .io_inputA              (pes_6_2_io_outputA[7:0]   ), //i
    .io_inputB              (pes_5_3_io_outputB[7:0]   ), //i
    .io_inputC              (pes_5_3_io_outputC[18:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_6_3), //i
    .io_outputA             (pes_6_3_io_outputA[7:0]   ), //o
    .io_outputB             (pes_6_3_io_outputB[7:0]   ), //o
    .io_outputC             (pes_6_3_io_outputC[18:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement_80 pes_6_4 (
    .io_inputA              (pes_6_3_io_outputA[7:0]   ), //i
    .io_inputB              (pes_5_4_io_outputB[7:0]   ), //i
    .io_inputC              (pes_5_4_io_outputC[18:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_6_4), //i
    .io_outputA             (pes_6_4_io_outputA[7:0]   ), //o
    .io_outputB             (pes_6_4_io_outputB[7:0]   ), //o
    .io_outputC             (pes_6_4_io_outputC[18:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement_80 pes_6_5 (
    .io_inputA              (pes_6_4_io_outputA[7:0]   ), //i
    .io_inputB              (pes_5_5_io_outputB[7:0]   ), //i
    .io_inputC              (pes_5_5_io_outputC[18:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_6_5), //i
    .io_outputA             (pes_6_5_io_outputA[7:0]   ), //o
    .io_outputB             (pes_6_5_io_outputB[7:0]   ), //o
    .io_outputC             (pes_6_5_io_outputC[18:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement_80 pes_6_6 (
    .io_inputA              (pes_6_5_io_outputA[7:0]   ), //i
    .io_inputB              (pes_5_6_io_outputB[7:0]   ), //i
    .io_inputC              (pes_5_6_io_outputC[18:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_6_6), //i
    .io_outputA             (pes_6_6_io_outputA[7:0]   ), //o
    .io_outputB             (pes_6_6_io_outputB[7:0]   ), //o
    .io_outputC             (pes_6_6_io_outputC[18:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement_80 pes_6_7 (
    .io_inputA              (pes_6_6_io_outputA[7:0]   ), //i
    .io_inputB              (pes_5_7_io_outputB[7:0]   ), //i
    .io_inputC              (pes_5_7_io_outputC[18:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_6_7), //i
    .io_outputA             (pes_6_7_io_outputA[7:0]   ), //o
    .io_outputB             (pes_6_7_io_outputB[7:0]   ), //o
    .io_outputC             (pes_6_7_io_outputC[18:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement_80 pes_6_8 (
    .io_inputA              (pes_6_7_io_outputA[7:0]   ), //i
    .io_inputB              (pes_5_8_io_outputB[7:0]   ), //i
    .io_inputC              (pes_5_8_io_outputC[18:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_6_8), //i
    .io_outputA             (pes_6_8_io_outputA[7:0]   ), //o
    .io_outputB             (pes_6_8_io_outputB[7:0]   ), //o
    .io_outputC             (pes_6_8_io_outputC[18:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement_80 pes_6_9 (
    .io_inputA              (pes_6_8_io_outputA[7:0]   ), //i
    .io_inputB              (pes_5_9_io_outputB[7:0]   ), //i
    .io_inputC              (pes_5_9_io_outputC[18:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_6_9), //i
    .io_outputA             (pes_6_9_io_outputA[7:0]   ), //o
    .io_outputB             (pes_6_9_io_outputB[7:0]   ), //o
    .io_outputC             (pes_6_9_io_outputC[18:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement_80 pes_6_10 (
    .io_inputA              (pes_6_9_io_outputA[7:0]    ), //i
    .io_inputB              (pes_5_10_io_outputB[7:0]   ), //i
    .io_inputC              (pes_5_10_io_outputC[18:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_6_10), //i
    .io_outputA             (pes_6_10_io_outputA[7:0]   ), //o
    .io_outputB             (pes_6_10_io_outputB[7:0]   ), //o
    .io_outputC             (pes_6_10_io_outputC[18:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_80 pes_6_11 (
    .io_inputA              (pes_6_10_io_outputA[7:0]   ), //i
    .io_inputB              (pes_5_11_io_outputB[7:0]   ), //i
    .io_inputC              (pes_5_11_io_outputC[18:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_6_11), //i
    .io_outputA             (pes_6_11_io_outputA[7:0]   ), //o
    .io_outputB             (pes_6_11_io_outputB[7:0]   ), //o
    .io_outputC             (pes_6_11_io_outputC[18:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_80 pes_6_12 (
    .io_inputA              (pes_6_11_io_outputA[7:0]   ), //i
    .io_inputB              (pes_5_12_io_outputB[7:0]   ), //i
    .io_inputC              (pes_5_12_io_outputC[18:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_6_12), //i
    .io_outputA             (pes_6_12_io_outputA[7:0]   ), //o
    .io_outputB             (pes_6_12_io_outputB[7:0]   ), //o
    .io_outputC             (pes_6_12_io_outputC[18:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_80 pes_6_13 (
    .io_inputA              (pes_6_12_io_outputA[7:0]   ), //i
    .io_inputB              (pes_5_13_io_outputB[7:0]   ), //i
    .io_inputC              (pes_5_13_io_outputC[18:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_6_13), //i
    .io_outputA             (pes_6_13_io_outputA[7:0]   ), //o
    .io_outputB             (pes_6_13_io_outputB[7:0]   ), //o
    .io_outputC             (pes_6_13_io_outputC[18:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_80 pes_6_14 (
    .io_inputA              (pes_6_13_io_outputA[7:0]   ), //i
    .io_inputB              (pes_5_14_io_outputB[7:0]   ), //i
    .io_inputC              (pes_5_14_io_outputC[18:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_6_14), //i
    .io_outputA             (pes_6_14_io_outputA[7:0]   ), //o
    .io_outputB             (pes_6_14_io_outputB[7:0]   ), //o
    .io_outputC             (pes_6_14_io_outputC[18:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_95 pes_6_15 (
    .io_inputA              (pes_6_14_io_outputA[7:0]   ), //i
    .io_inputB              (pes_5_15_io_outputB[7:0]   ), //i
    .io_inputC              (pes_5_15_io_outputC[18:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_6_15), //i
    .io_outputB             (pes_6_15_io_outputB[7:0]   ), //o
    .io_outputC             (pes_6_15_io_outputC[18:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_80 pes_7_0 (
    .io_inputA              (skewBuffer_io_output_7[7:0]), //i
    .io_inputB              (pes_6_0_io_outputB[7:0]    ), //i
    .io_inputC              (pes_6_0_io_outputC[18:0]   ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_7_0 ), //i
    .io_outputA             (pes_7_0_io_outputA[7:0]    ), //o
    .io_outputB             (pes_7_0_io_outputB[7:0]    ), //o
    .io_outputC             (pes_7_0_io_outputC[18:0]   ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_80 pes_7_1 (
    .io_inputA              (pes_7_0_io_outputA[7:0]   ), //i
    .io_inputB              (pes_6_1_io_outputB[7:0]   ), //i
    .io_inputC              (pes_6_1_io_outputC[18:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_7_1), //i
    .io_outputA             (pes_7_1_io_outputA[7:0]   ), //o
    .io_outputB             (pes_7_1_io_outputB[7:0]   ), //o
    .io_outputC             (pes_7_1_io_outputC[18:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement_80 pes_7_2 (
    .io_inputA              (pes_7_1_io_outputA[7:0]   ), //i
    .io_inputB              (pes_6_2_io_outputB[7:0]   ), //i
    .io_inputC              (pes_6_2_io_outputC[18:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_7_2), //i
    .io_outputA             (pes_7_2_io_outputA[7:0]   ), //o
    .io_outputB             (pes_7_2_io_outputB[7:0]   ), //o
    .io_outputC             (pes_7_2_io_outputC[18:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement_80 pes_7_3 (
    .io_inputA              (pes_7_2_io_outputA[7:0]   ), //i
    .io_inputB              (pes_6_3_io_outputB[7:0]   ), //i
    .io_inputC              (pes_6_3_io_outputC[18:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_7_3), //i
    .io_outputA             (pes_7_3_io_outputA[7:0]   ), //o
    .io_outputB             (pes_7_3_io_outputB[7:0]   ), //o
    .io_outputC             (pes_7_3_io_outputC[18:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement_80 pes_7_4 (
    .io_inputA              (pes_7_3_io_outputA[7:0]   ), //i
    .io_inputB              (pes_6_4_io_outputB[7:0]   ), //i
    .io_inputC              (pes_6_4_io_outputC[18:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_7_4), //i
    .io_outputA             (pes_7_4_io_outputA[7:0]   ), //o
    .io_outputB             (pes_7_4_io_outputB[7:0]   ), //o
    .io_outputC             (pes_7_4_io_outputC[18:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement_80 pes_7_5 (
    .io_inputA              (pes_7_4_io_outputA[7:0]   ), //i
    .io_inputB              (pes_6_5_io_outputB[7:0]   ), //i
    .io_inputC              (pes_6_5_io_outputC[18:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_7_5), //i
    .io_outputA             (pes_7_5_io_outputA[7:0]   ), //o
    .io_outputB             (pes_7_5_io_outputB[7:0]   ), //o
    .io_outputC             (pes_7_5_io_outputC[18:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement_80 pes_7_6 (
    .io_inputA              (pes_7_5_io_outputA[7:0]   ), //i
    .io_inputB              (pes_6_6_io_outputB[7:0]   ), //i
    .io_inputC              (pes_6_6_io_outputC[18:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_7_6), //i
    .io_outputA             (pes_7_6_io_outputA[7:0]   ), //o
    .io_outputB             (pes_7_6_io_outputB[7:0]   ), //o
    .io_outputC             (pes_7_6_io_outputC[18:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement_80 pes_7_7 (
    .io_inputA              (pes_7_6_io_outputA[7:0]   ), //i
    .io_inputB              (pes_6_7_io_outputB[7:0]   ), //i
    .io_inputC              (pes_6_7_io_outputC[18:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_7_7), //i
    .io_outputA             (pes_7_7_io_outputA[7:0]   ), //o
    .io_outputB             (pes_7_7_io_outputB[7:0]   ), //o
    .io_outputC             (pes_7_7_io_outputC[18:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement_80 pes_7_8 (
    .io_inputA              (pes_7_7_io_outputA[7:0]   ), //i
    .io_inputB              (pes_6_8_io_outputB[7:0]   ), //i
    .io_inputC              (pes_6_8_io_outputC[18:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_7_8), //i
    .io_outputA             (pes_7_8_io_outputA[7:0]   ), //o
    .io_outputB             (pes_7_8_io_outputB[7:0]   ), //o
    .io_outputC             (pes_7_8_io_outputC[18:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement_80 pes_7_9 (
    .io_inputA              (pes_7_8_io_outputA[7:0]   ), //i
    .io_inputB              (pes_6_9_io_outputB[7:0]   ), //i
    .io_inputC              (pes_6_9_io_outputC[18:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_7_9), //i
    .io_outputA             (pes_7_9_io_outputA[7:0]   ), //o
    .io_outputB             (pes_7_9_io_outputB[7:0]   ), //o
    .io_outputC             (pes_7_9_io_outputC[18:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement_80 pes_7_10 (
    .io_inputA              (pes_7_9_io_outputA[7:0]    ), //i
    .io_inputB              (pes_6_10_io_outputB[7:0]   ), //i
    .io_inputC              (pes_6_10_io_outputC[18:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_7_10), //i
    .io_outputA             (pes_7_10_io_outputA[7:0]   ), //o
    .io_outputB             (pes_7_10_io_outputB[7:0]   ), //o
    .io_outputC             (pes_7_10_io_outputC[18:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_80 pes_7_11 (
    .io_inputA              (pes_7_10_io_outputA[7:0]   ), //i
    .io_inputB              (pes_6_11_io_outputB[7:0]   ), //i
    .io_inputC              (pes_6_11_io_outputC[18:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_7_11), //i
    .io_outputA             (pes_7_11_io_outputA[7:0]   ), //o
    .io_outputB             (pes_7_11_io_outputB[7:0]   ), //o
    .io_outputC             (pes_7_11_io_outputC[18:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_80 pes_7_12 (
    .io_inputA              (pes_7_11_io_outputA[7:0]   ), //i
    .io_inputB              (pes_6_12_io_outputB[7:0]   ), //i
    .io_inputC              (pes_6_12_io_outputC[18:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_7_12), //i
    .io_outputA             (pes_7_12_io_outputA[7:0]   ), //o
    .io_outputB             (pes_7_12_io_outputB[7:0]   ), //o
    .io_outputC             (pes_7_12_io_outputC[18:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_80 pes_7_13 (
    .io_inputA              (pes_7_12_io_outputA[7:0]   ), //i
    .io_inputB              (pes_6_13_io_outputB[7:0]   ), //i
    .io_inputC              (pes_6_13_io_outputC[18:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_7_13), //i
    .io_outputA             (pes_7_13_io_outputA[7:0]   ), //o
    .io_outputB             (pes_7_13_io_outputB[7:0]   ), //o
    .io_outputC             (pes_7_13_io_outputC[18:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_80 pes_7_14 (
    .io_inputA              (pes_7_13_io_outputA[7:0]   ), //i
    .io_inputB              (pes_6_14_io_outputB[7:0]   ), //i
    .io_inputC              (pes_6_14_io_outputC[18:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_7_14), //i
    .io_outputA             (pes_7_14_io_outputA[7:0]   ), //o
    .io_outputB             (pes_7_14_io_outputB[7:0]   ), //o
    .io_outputC             (pes_7_14_io_outputC[18:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_95 pes_7_15 (
    .io_inputA              (pes_7_14_io_outputA[7:0]   ), //i
    .io_inputB              (pes_6_15_io_outputB[7:0]   ), //i
    .io_inputC              (pes_6_15_io_outputC[18:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_7_15), //i
    .io_outputB             (pes_7_15_io_outputB[7:0]   ), //o
    .io_outputC             (pes_7_15_io_outputC[18:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_128 pes_8_0 (
    .io_inputA              (skewBuffer_io_output_8[7:0]), //i
    .io_inputB              (pes_7_0_io_outputB[7:0]    ), //i
    .io_inputC              (pes_7_0_io_outputC[18:0]   ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_8_0 ), //i
    .io_outputA             (pes_8_0_io_outputA[7:0]    ), //o
    .io_outputB             (pes_8_0_io_outputB[7:0]    ), //o
    .io_outputC             (pes_8_0_io_outputC[19:0]   ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_128 pes_8_1 (
    .io_inputA              (pes_8_0_io_outputA[7:0]   ), //i
    .io_inputB              (pes_7_1_io_outputB[7:0]   ), //i
    .io_inputC              (pes_7_1_io_outputC[18:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_8_1), //i
    .io_outputA             (pes_8_1_io_outputA[7:0]   ), //o
    .io_outputB             (pes_8_1_io_outputB[7:0]   ), //o
    .io_outputC             (pes_8_1_io_outputC[19:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement_128 pes_8_2 (
    .io_inputA              (pes_8_1_io_outputA[7:0]   ), //i
    .io_inputB              (pes_7_2_io_outputB[7:0]   ), //i
    .io_inputC              (pes_7_2_io_outputC[18:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_8_2), //i
    .io_outputA             (pes_8_2_io_outputA[7:0]   ), //o
    .io_outputB             (pes_8_2_io_outputB[7:0]   ), //o
    .io_outputC             (pes_8_2_io_outputC[19:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement_128 pes_8_3 (
    .io_inputA              (pes_8_2_io_outputA[7:0]   ), //i
    .io_inputB              (pes_7_3_io_outputB[7:0]   ), //i
    .io_inputC              (pes_7_3_io_outputC[18:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_8_3), //i
    .io_outputA             (pes_8_3_io_outputA[7:0]   ), //o
    .io_outputB             (pes_8_3_io_outputB[7:0]   ), //o
    .io_outputC             (pes_8_3_io_outputC[19:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement_128 pes_8_4 (
    .io_inputA              (pes_8_3_io_outputA[7:0]   ), //i
    .io_inputB              (pes_7_4_io_outputB[7:0]   ), //i
    .io_inputC              (pes_7_4_io_outputC[18:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_8_4), //i
    .io_outputA             (pes_8_4_io_outputA[7:0]   ), //o
    .io_outputB             (pes_8_4_io_outputB[7:0]   ), //o
    .io_outputC             (pes_8_4_io_outputC[19:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement_128 pes_8_5 (
    .io_inputA              (pes_8_4_io_outputA[7:0]   ), //i
    .io_inputB              (pes_7_5_io_outputB[7:0]   ), //i
    .io_inputC              (pes_7_5_io_outputC[18:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_8_5), //i
    .io_outputA             (pes_8_5_io_outputA[7:0]   ), //o
    .io_outputB             (pes_8_5_io_outputB[7:0]   ), //o
    .io_outputC             (pes_8_5_io_outputC[19:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement_128 pes_8_6 (
    .io_inputA              (pes_8_5_io_outputA[7:0]   ), //i
    .io_inputB              (pes_7_6_io_outputB[7:0]   ), //i
    .io_inputC              (pes_7_6_io_outputC[18:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_8_6), //i
    .io_outputA             (pes_8_6_io_outputA[7:0]   ), //o
    .io_outputB             (pes_8_6_io_outputB[7:0]   ), //o
    .io_outputC             (pes_8_6_io_outputC[19:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement_128 pes_8_7 (
    .io_inputA              (pes_8_6_io_outputA[7:0]   ), //i
    .io_inputB              (pes_7_7_io_outputB[7:0]   ), //i
    .io_inputC              (pes_7_7_io_outputC[18:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_8_7), //i
    .io_outputA             (pes_8_7_io_outputA[7:0]   ), //o
    .io_outputB             (pes_8_7_io_outputB[7:0]   ), //o
    .io_outputC             (pes_8_7_io_outputC[19:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement_128 pes_8_8 (
    .io_inputA              (pes_8_7_io_outputA[7:0]   ), //i
    .io_inputB              (pes_7_8_io_outputB[7:0]   ), //i
    .io_inputC              (pes_7_8_io_outputC[18:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_8_8), //i
    .io_outputA             (pes_8_8_io_outputA[7:0]   ), //o
    .io_outputB             (pes_8_8_io_outputB[7:0]   ), //o
    .io_outputC             (pes_8_8_io_outputC[19:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement_128 pes_8_9 (
    .io_inputA              (pes_8_8_io_outputA[7:0]   ), //i
    .io_inputB              (pes_7_9_io_outputB[7:0]   ), //i
    .io_inputC              (pes_7_9_io_outputC[18:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_8_9), //i
    .io_outputA             (pes_8_9_io_outputA[7:0]   ), //o
    .io_outputB             (pes_8_9_io_outputB[7:0]   ), //o
    .io_outputC             (pes_8_9_io_outputC[19:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement_128 pes_8_10 (
    .io_inputA              (pes_8_9_io_outputA[7:0]    ), //i
    .io_inputB              (pes_7_10_io_outputB[7:0]   ), //i
    .io_inputC              (pes_7_10_io_outputC[18:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_8_10), //i
    .io_outputA             (pes_8_10_io_outputA[7:0]   ), //o
    .io_outputB             (pes_8_10_io_outputB[7:0]   ), //o
    .io_outputC             (pes_8_10_io_outputC[19:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_128 pes_8_11 (
    .io_inputA              (pes_8_10_io_outputA[7:0]   ), //i
    .io_inputB              (pes_7_11_io_outputB[7:0]   ), //i
    .io_inputC              (pes_7_11_io_outputC[18:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_8_11), //i
    .io_outputA             (pes_8_11_io_outputA[7:0]   ), //o
    .io_outputB             (pes_8_11_io_outputB[7:0]   ), //o
    .io_outputC             (pes_8_11_io_outputC[19:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_128 pes_8_12 (
    .io_inputA              (pes_8_11_io_outputA[7:0]   ), //i
    .io_inputB              (pes_7_12_io_outputB[7:0]   ), //i
    .io_inputC              (pes_7_12_io_outputC[18:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_8_12), //i
    .io_outputA             (pes_8_12_io_outputA[7:0]   ), //o
    .io_outputB             (pes_8_12_io_outputB[7:0]   ), //o
    .io_outputC             (pes_8_12_io_outputC[19:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_128 pes_8_13 (
    .io_inputA              (pes_8_12_io_outputA[7:0]   ), //i
    .io_inputB              (pes_7_13_io_outputB[7:0]   ), //i
    .io_inputC              (pes_7_13_io_outputC[18:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_8_13), //i
    .io_outputA             (pes_8_13_io_outputA[7:0]   ), //o
    .io_outputB             (pes_8_13_io_outputB[7:0]   ), //o
    .io_outputC             (pes_8_13_io_outputC[19:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_128 pes_8_14 (
    .io_inputA              (pes_8_13_io_outputA[7:0]   ), //i
    .io_inputB              (pes_7_14_io_outputB[7:0]   ), //i
    .io_inputC              (pes_7_14_io_outputC[18:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_8_14), //i
    .io_outputA             (pes_8_14_io_outputA[7:0]   ), //o
    .io_outputB             (pes_8_14_io_outputB[7:0]   ), //o
    .io_outputC             (pes_8_14_io_outputC[19:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_143 pes_8_15 (
    .io_inputA              (pes_8_14_io_outputA[7:0]   ), //i
    .io_inputB              (pes_7_15_io_outputB[7:0]   ), //i
    .io_inputC              (pes_7_15_io_outputC[18:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_8_15), //i
    .io_outputB             (pes_8_15_io_outputB[7:0]   ), //o
    .io_outputC             (pes_8_15_io_outputC[19:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_144 pes_9_0 (
    .io_inputA              (skewBuffer_io_output_9[7:0]), //i
    .io_inputB              (pes_8_0_io_outputB[7:0]    ), //i
    .io_inputC              (pes_8_0_io_outputC[19:0]   ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_9_0 ), //i
    .io_outputA             (pes_9_0_io_outputA[7:0]    ), //o
    .io_outputB             (pes_9_0_io_outputB[7:0]    ), //o
    .io_outputC             (pes_9_0_io_outputC[19:0]   ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_144 pes_9_1 (
    .io_inputA              (pes_9_0_io_outputA[7:0]   ), //i
    .io_inputB              (pes_8_1_io_outputB[7:0]   ), //i
    .io_inputC              (pes_8_1_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_9_1), //i
    .io_outputA             (pes_9_1_io_outputA[7:0]   ), //o
    .io_outputB             (pes_9_1_io_outputB[7:0]   ), //o
    .io_outputC             (pes_9_1_io_outputC[19:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement_144 pes_9_2 (
    .io_inputA              (pes_9_1_io_outputA[7:0]   ), //i
    .io_inputB              (pes_8_2_io_outputB[7:0]   ), //i
    .io_inputC              (pes_8_2_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_9_2), //i
    .io_outputA             (pes_9_2_io_outputA[7:0]   ), //o
    .io_outputB             (pes_9_2_io_outputB[7:0]   ), //o
    .io_outputC             (pes_9_2_io_outputC[19:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement_144 pes_9_3 (
    .io_inputA              (pes_9_2_io_outputA[7:0]   ), //i
    .io_inputB              (pes_8_3_io_outputB[7:0]   ), //i
    .io_inputC              (pes_8_3_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_9_3), //i
    .io_outputA             (pes_9_3_io_outputA[7:0]   ), //o
    .io_outputB             (pes_9_3_io_outputB[7:0]   ), //o
    .io_outputC             (pes_9_3_io_outputC[19:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement_144 pes_9_4 (
    .io_inputA              (pes_9_3_io_outputA[7:0]   ), //i
    .io_inputB              (pes_8_4_io_outputB[7:0]   ), //i
    .io_inputC              (pes_8_4_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_9_4), //i
    .io_outputA             (pes_9_4_io_outputA[7:0]   ), //o
    .io_outputB             (pes_9_4_io_outputB[7:0]   ), //o
    .io_outputC             (pes_9_4_io_outputC[19:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement_144 pes_9_5 (
    .io_inputA              (pes_9_4_io_outputA[7:0]   ), //i
    .io_inputB              (pes_8_5_io_outputB[7:0]   ), //i
    .io_inputC              (pes_8_5_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_9_5), //i
    .io_outputA             (pes_9_5_io_outputA[7:0]   ), //o
    .io_outputB             (pes_9_5_io_outputB[7:0]   ), //o
    .io_outputC             (pes_9_5_io_outputC[19:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement_144 pes_9_6 (
    .io_inputA              (pes_9_5_io_outputA[7:0]   ), //i
    .io_inputB              (pes_8_6_io_outputB[7:0]   ), //i
    .io_inputC              (pes_8_6_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_9_6), //i
    .io_outputA             (pes_9_6_io_outputA[7:0]   ), //o
    .io_outputB             (pes_9_6_io_outputB[7:0]   ), //o
    .io_outputC             (pes_9_6_io_outputC[19:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement_144 pes_9_7 (
    .io_inputA              (pes_9_6_io_outputA[7:0]   ), //i
    .io_inputB              (pes_8_7_io_outputB[7:0]   ), //i
    .io_inputC              (pes_8_7_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_9_7), //i
    .io_outputA             (pes_9_7_io_outputA[7:0]   ), //o
    .io_outputB             (pes_9_7_io_outputB[7:0]   ), //o
    .io_outputC             (pes_9_7_io_outputC[19:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement_144 pes_9_8 (
    .io_inputA              (pes_9_7_io_outputA[7:0]   ), //i
    .io_inputB              (pes_8_8_io_outputB[7:0]   ), //i
    .io_inputC              (pes_8_8_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_9_8), //i
    .io_outputA             (pes_9_8_io_outputA[7:0]   ), //o
    .io_outputB             (pes_9_8_io_outputB[7:0]   ), //o
    .io_outputC             (pes_9_8_io_outputC[19:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement_144 pes_9_9 (
    .io_inputA              (pes_9_8_io_outputA[7:0]   ), //i
    .io_inputB              (pes_8_9_io_outputB[7:0]   ), //i
    .io_inputC              (pes_8_9_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_9_9), //i
    .io_outputA             (pes_9_9_io_outputA[7:0]   ), //o
    .io_outputB             (pes_9_9_io_outputB[7:0]   ), //o
    .io_outputC             (pes_9_9_io_outputC[19:0]  ), //o
    .clk                    (clk                       ), //i
    .reset                  (reset                     )  //i
  );
  ProcessingElement_144 pes_9_10 (
    .io_inputA              (pes_9_9_io_outputA[7:0]    ), //i
    .io_inputB              (pes_8_10_io_outputB[7:0]   ), //i
    .io_inputC              (pes_8_10_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_9_10), //i
    .io_outputA             (pes_9_10_io_outputA[7:0]   ), //o
    .io_outputB             (pes_9_10_io_outputB[7:0]   ), //o
    .io_outputC             (pes_9_10_io_outputC[19:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_144 pes_9_11 (
    .io_inputA              (pes_9_10_io_outputA[7:0]   ), //i
    .io_inputB              (pes_8_11_io_outputB[7:0]   ), //i
    .io_inputC              (pes_8_11_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_9_11), //i
    .io_outputA             (pes_9_11_io_outputA[7:0]   ), //o
    .io_outputB             (pes_9_11_io_outputB[7:0]   ), //o
    .io_outputC             (pes_9_11_io_outputC[19:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_144 pes_9_12 (
    .io_inputA              (pes_9_11_io_outputA[7:0]   ), //i
    .io_inputB              (pes_8_12_io_outputB[7:0]   ), //i
    .io_inputC              (pes_8_12_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_9_12), //i
    .io_outputA             (pes_9_12_io_outputA[7:0]   ), //o
    .io_outputB             (pes_9_12_io_outputB[7:0]   ), //o
    .io_outputC             (pes_9_12_io_outputC[19:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_144 pes_9_13 (
    .io_inputA              (pes_9_12_io_outputA[7:0]   ), //i
    .io_inputB              (pes_8_13_io_outputB[7:0]   ), //i
    .io_inputC              (pes_8_13_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_9_13), //i
    .io_outputA             (pes_9_13_io_outputA[7:0]   ), //o
    .io_outputB             (pes_9_13_io_outputB[7:0]   ), //o
    .io_outputC             (pes_9_13_io_outputC[19:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_144 pes_9_14 (
    .io_inputA              (pes_9_13_io_outputA[7:0]   ), //i
    .io_inputB              (pes_8_14_io_outputB[7:0]   ), //i
    .io_inputC              (pes_8_14_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_9_14), //i
    .io_outputA             (pes_9_14_io_outputA[7:0]   ), //o
    .io_outputB             (pes_9_14_io_outputB[7:0]   ), //o
    .io_outputC             (pes_9_14_io_outputC[19:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_159 pes_9_15 (
    .io_inputA              (pes_9_14_io_outputA[7:0]   ), //i
    .io_inputB              (pes_8_15_io_outputB[7:0]   ), //i
    .io_inputC              (pes_8_15_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_9_15), //i
    .io_outputB             (pes_9_15_io_outputB[7:0]   ), //o
    .io_outputC             (pes_9_15_io_outputC[19:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_144 pes_10_0 (
    .io_inputA              (skewBuffer_io_output_10[7:0]), //i
    .io_inputB              (pes_9_0_io_outputB[7:0]     ), //i
    .io_inputC              (pes_9_0_io_outputC[19:0]    ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_10_0 ), //i
    .io_outputA             (pes_10_0_io_outputA[7:0]    ), //o
    .io_outputB             (pes_10_0_io_outputB[7:0]    ), //o
    .io_outputC             (pes_10_0_io_outputC[19:0]   ), //o
    .clk                    (clk                         ), //i
    .reset                  (reset                       )  //i
  );
  ProcessingElement_144 pes_10_1 (
    .io_inputA              (pes_10_0_io_outputA[7:0]   ), //i
    .io_inputB              (pes_9_1_io_outputB[7:0]    ), //i
    .io_inputC              (pes_9_1_io_outputC[19:0]   ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_10_1), //i
    .io_outputA             (pes_10_1_io_outputA[7:0]   ), //o
    .io_outputB             (pes_10_1_io_outputB[7:0]   ), //o
    .io_outputC             (pes_10_1_io_outputC[19:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_144 pes_10_2 (
    .io_inputA              (pes_10_1_io_outputA[7:0]   ), //i
    .io_inputB              (pes_9_2_io_outputB[7:0]    ), //i
    .io_inputC              (pes_9_2_io_outputC[19:0]   ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_10_2), //i
    .io_outputA             (pes_10_2_io_outputA[7:0]   ), //o
    .io_outputB             (pes_10_2_io_outputB[7:0]   ), //o
    .io_outputC             (pes_10_2_io_outputC[19:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_144 pes_10_3 (
    .io_inputA              (pes_10_2_io_outputA[7:0]   ), //i
    .io_inputB              (pes_9_3_io_outputB[7:0]    ), //i
    .io_inputC              (pes_9_3_io_outputC[19:0]   ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_10_3), //i
    .io_outputA             (pes_10_3_io_outputA[7:0]   ), //o
    .io_outputB             (pes_10_3_io_outputB[7:0]   ), //o
    .io_outputC             (pes_10_3_io_outputC[19:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_144 pes_10_4 (
    .io_inputA              (pes_10_3_io_outputA[7:0]   ), //i
    .io_inputB              (pes_9_4_io_outputB[7:0]    ), //i
    .io_inputC              (pes_9_4_io_outputC[19:0]   ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_10_4), //i
    .io_outputA             (pes_10_4_io_outputA[7:0]   ), //o
    .io_outputB             (pes_10_4_io_outputB[7:0]   ), //o
    .io_outputC             (pes_10_4_io_outputC[19:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_144 pes_10_5 (
    .io_inputA              (pes_10_4_io_outputA[7:0]   ), //i
    .io_inputB              (pes_9_5_io_outputB[7:0]    ), //i
    .io_inputC              (pes_9_5_io_outputC[19:0]   ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_10_5), //i
    .io_outputA             (pes_10_5_io_outputA[7:0]   ), //o
    .io_outputB             (pes_10_5_io_outputB[7:0]   ), //o
    .io_outputC             (pes_10_5_io_outputC[19:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_144 pes_10_6 (
    .io_inputA              (pes_10_5_io_outputA[7:0]   ), //i
    .io_inputB              (pes_9_6_io_outputB[7:0]    ), //i
    .io_inputC              (pes_9_6_io_outputC[19:0]   ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_10_6), //i
    .io_outputA             (pes_10_6_io_outputA[7:0]   ), //o
    .io_outputB             (pes_10_6_io_outputB[7:0]   ), //o
    .io_outputC             (pes_10_6_io_outputC[19:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_144 pes_10_7 (
    .io_inputA              (pes_10_6_io_outputA[7:0]   ), //i
    .io_inputB              (pes_9_7_io_outputB[7:0]    ), //i
    .io_inputC              (pes_9_7_io_outputC[19:0]   ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_10_7), //i
    .io_outputA             (pes_10_7_io_outputA[7:0]   ), //o
    .io_outputB             (pes_10_7_io_outputB[7:0]   ), //o
    .io_outputC             (pes_10_7_io_outputC[19:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_144 pes_10_8 (
    .io_inputA              (pes_10_7_io_outputA[7:0]   ), //i
    .io_inputB              (pes_9_8_io_outputB[7:0]    ), //i
    .io_inputC              (pes_9_8_io_outputC[19:0]   ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_10_8), //i
    .io_outputA             (pes_10_8_io_outputA[7:0]   ), //o
    .io_outputB             (pes_10_8_io_outputB[7:0]   ), //o
    .io_outputC             (pes_10_8_io_outputC[19:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_144 pes_10_9 (
    .io_inputA              (pes_10_8_io_outputA[7:0]   ), //i
    .io_inputB              (pes_9_9_io_outputB[7:0]    ), //i
    .io_inputC              (pes_9_9_io_outputC[19:0]   ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_10_9), //i
    .io_outputA             (pes_10_9_io_outputA[7:0]   ), //o
    .io_outputB             (pes_10_9_io_outputB[7:0]   ), //o
    .io_outputC             (pes_10_9_io_outputC[19:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_144 pes_10_10 (
    .io_inputA              (pes_10_9_io_outputA[7:0]    ), //i
    .io_inputB              (pes_9_10_io_outputB[7:0]    ), //i
    .io_inputC              (pes_9_10_io_outputC[19:0]   ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_10_10), //i
    .io_outputA             (pes_10_10_io_outputA[7:0]   ), //o
    .io_outputB             (pes_10_10_io_outputB[7:0]   ), //o
    .io_outputC             (pes_10_10_io_outputC[19:0]  ), //o
    .clk                    (clk                         ), //i
    .reset                  (reset                       )  //i
  );
  ProcessingElement_144 pes_10_11 (
    .io_inputA              (pes_10_10_io_outputA[7:0]   ), //i
    .io_inputB              (pes_9_11_io_outputB[7:0]    ), //i
    .io_inputC              (pes_9_11_io_outputC[19:0]   ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_10_11), //i
    .io_outputA             (pes_10_11_io_outputA[7:0]   ), //o
    .io_outputB             (pes_10_11_io_outputB[7:0]   ), //o
    .io_outputC             (pes_10_11_io_outputC[19:0]  ), //o
    .clk                    (clk                         ), //i
    .reset                  (reset                       )  //i
  );
  ProcessingElement_144 pes_10_12 (
    .io_inputA              (pes_10_11_io_outputA[7:0]   ), //i
    .io_inputB              (pes_9_12_io_outputB[7:0]    ), //i
    .io_inputC              (pes_9_12_io_outputC[19:0]   ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_10_12), //i
    .io_outputA             (pes_10_12_io_outputA[7:0]   ), //o
    .io_outputB             (pes_10_12_io_outputB[7:0]   ), //o
    .io_outputC             (pes_10_12_io_outputC[19:0]  ), //o
    .clk                    (clk                         ), //i
    .reset                  (reset                       )  //i
  );
  ProcessingElement_144 pes_10_13 (
    .io_inputA              (pes_10_12_io_outputA[7:0]   ), //i
    .io_inputB              (pes_9_13_io_outputB[7:0]    ), //i
    .io_inputC              (pes_9_13_io_outputC[19:0]   ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_10_13), //i
    .io_outputA             (pes_10_13_io_outputA[7:0]   ), //o
    .io_outputB             (pes_10_13_io_outputB[7:0]   ), //o
    .io_outputC             (pes_10_13_io_outputC[19:0]  ), //o
    .clk                    (clk                         ), //i
    .reset                  (reset                       )  //i
  );
  ProcessingElement_144 pes_10_14 (
    .io_inputA              (pes_10_13_io_outputA[7:0]   ), //i
    .io_inputB              (pes_9_14_io_outputB[7:0]    ), //i
    .io_inputC              (pes_9_14_io_outputC[19:0]   ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_10_14), //i
    .io_outputA             (pes_10_14_io_outputA[7:0]   ), //o
    .io_outputB             (pes_10_14_io_outputB[7:0]   ), //o
    .io_outputC             (pes_10_14_io_outputC[19:0]  ), //o
    .clk                    (clk                         ), //i
    .reset                  (reset                       )  //i
  );
  ProcessingElement_159 pes_10_15 (
    .io_inputA              (pes_10_14_io_outputA[7:0]   ), //i
    .io_inputB              (pes_9_15_io_outputB[7:0]    ), //i
    .io_inputC              (pes_9_15_io_outputC[19:0]   ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_10_15), //i
    .io_outputB             (pes_10_15_io_outputB[7:0]   ), //o
    .io_outputC             (pes_10_15_io_outputC[19:0]  ), //o
    .clk                    (clk                         ), //i
    .reset                  (reset                       )  //i
  );
  ProcessingElement_144 pes_11_0 (
    .io_inputA              (skewBuffer_io_output_11[7:0]), //i
    .io_inputB              (pes_10_0_io_outputB[7:0]    ), //i
    .io_inputC              (pes_10_0_io_outputC[19:0]   ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_11_0 ), //i
    .io_outputA             (pes_11_0_io_outputA[7:0]    ), //o
    .io_outputB             (pes_11_0_io_outputB[7:0]    ), //o
    .io_outputC             (pes_11_0_io_outputC[19:0]   ), //o
    .clk                    (clk                         ), //i
    .reset                  (reset                       )  //i
  );
  ProcessingElement_144 pes_11_1 (
    .io_inputA              (pes_11_0_io_outputA[7:0]   ), //i
    .io_inputB              (pes_10_1_io_outputB[7:0]   ), //i
    .io_inputC              (pes_10_1_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_11_1), //i
    .io_outputA             (pes_11_1_io_outputA[7:0]   ), //o
    .io_outputB             (pes_11_1_io_outputB[7:0]   ), //o
    .io_outputC             (pes_11_1_io_outputC[19:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_144 pes_11_2 (
    .io_inputA              (pes_11_1_io_outputA[7:0]   ), //i
    .io_inputB              (pes_10_2_io_outputB[7:0]   ), //i
    .io_inputC              (pes_10_2_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_11_2), //i
    .io_outputA             (pes_11_2_io_outputA[7:0]   ), //o
    .io_outputB             (pes_11_2_io_outputB[7:0]   ), //o
    .io_outputC             (pes_11_2_io_outputC[19:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_144 pes_11_3 (
    .io_inputA              (pes_11_2_io_outputA[7:0]   ), //i
    .io_inputB              (pes_10_3_io_outputB[7:0]   ), //i
    .io_inputC              (pes_10_3_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_11_3), //i
    .io_outputA             (pes_11_3_io_outputA[7:0]   ), //o
    .io_outputB             (pes_11_3_io_outputB[7:0]   ), //o
    .io_outputC             (pes_11_3_io_outputC[19:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_144 pes_11_4 (
    .io_inputA              (pes_11_3_io_outputA[7:0]   ), //i
    .io_inputB              (pes_10_4_io_outputB[7:0]   ), //i
    .io_inputC              (pes_10_4_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_11_4), //i
    .io_outputA             (pes_11_4_io_outputA[7:0]   ), //o
    .io_outputB             (pes_11_4_io_outputB[7:0]   ), //o
    .io_outputC             (pes_11_4_io_outputC[19:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_144 pes_11_5 (
    .io_inputA              (pes_11_4_io_outputA[7:0]   ), //i
    .io_inputB              (pes_10_5_io_outputB[7:0]   ), //i
    .io_inputC              (pes_10_5_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_11_5), //i
    .io_outputA             (pes_11_5_io_outputA[7:0]   ), //o
    .io_outputB             (pes_11_5_io_outputB[7:0]   ), //o
    .io_outputC             (pes_11_5_io_outputC[19:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_144 pes_11_6 (
    .io_inputA              (pes_11_5_io_outputA[7:0]   ), //i
    .io_inputB              (pes_10_6_io_outputB[7:0]   ), //i
    .io_inputC              (pes_10_6_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_11_6), //i
    .io_outputA             (pes_11_6_io_outputA[7:0]   ), //o
    .io_outputB             (pes_11_6_io_outputB[7:0]   ), //o
    .io_outputC             (pes_11_6_io_outputC[19:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_144 pes_11_7 (
    .io_inputA              (pes_11_6_io_outputA[7:0]   ), //i
    .io_inputB              (pes_10_7_io_outputB[7:0]   ), //i
    .io_inputC              (pes_10_7_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_11_7), //i
    .io_outputA             (pes_11_7_io_outputA[7:0]   ), //o
    .io_outputB             (pes_11_7_io_outputB[7:0]   ), //o
    .io_outputC             (pes_11_7_io_outputC[19:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_144 pes_11_8 (
    .io_inputA              (pes_11_7_io_outputA[7:0]   ), //i
    .io_inputB              (pes_10_8_io_outputB[7:0]   ), //i
    .io_inputC              (pes_10_8_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_11_8), //i
    .io_outputA             (pes_11_8_io_outputA[7:0]   ), //o
    .io_outputB             (pes_11_8_io_outputB[7:0]   ), //o
    .io_outputC             (pes_11_8_io_outputC[19:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_144 pes_11_9 (
    .io_inputA              (pes_11_8_io_outputA[7:0]   ), //i
    .io_inputB              (pes_10_9_io_outputB[7:0]   ), //i
    .io_inputC              (pes_10_9_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_11_9), //i
    .io_outputA             (pes_11_9_io_outputA[7:0]   ), //o
    .io_outputB             (pes_11_9_io_outputB[7:0]   ), //o
    .io_outputC             (pes_11_9_io_outputC[19:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_144 pes_11_10 (
    .io_inputA              (pes_11_9_io_outputA[7:0]    ), //i
    .io_inputB              (pes_10_10_io_outputB[7:0]   ), //i
    .io_inputC              (pes_10_10_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_11_10), //i
    .io_outputA             (pes_11_10_io_outputA[7:0]   ), //o
    .io_outputB             (pes_11_10_io_outputB[7:0]   ), //o
    .io_outputC             (pes_11_10_io_outputC[19:0]  ), //o
    .clk                    (clk                         ), //i
    .reset                  (reset                       )  //i
  );
  ProcessingElement_144 pes_11_11 (
    .io_inputA              (pes_11_10_io_outputA[7:0]   ), //i
    .io_inputB              (pes_10_11_io_outputB[7:0]   ), //i
    .io_inputC              (pes_10_11_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_11_11), //i
    .io_outputA             (pes_11_11_io_outputA[7:0]   ), //o
    .io_outputB             (pes_11_11_io_outputB[7:0]   ), //o
    .io_outputC             (pes_11_11_io_outputC[19:0]  ), //o
    .clk                    (clk                         ), //i
    .reset                  (reset                       )  //i
  );
  ProcessingElement_144 pes_11_12 (
    .io_inputA              (pes_11_11_io_outputA[7:0]   ), //i
    .io_inputB              (pes_10_12_io_outputB[7:0]   ), //i
    .io_inputC              (pes_10_12_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_11_12), //i
    .io_outputA             (pes_11_12_io_outputA[7:0]   ), //o
    .io_outputB             (pes_11_12_io_outputB[7:0]   ), //o
    .io_outputC             (pes_11_12_io_outputC[19:0]  ), //o
    .clk                    (clk                         ), //i
    .reset                  (reset                       )  //i
  );
  ProcessingElement_144 pes_11_13 (
    .io_inputA              (pes_11_12_io_outputA[7:0]   ), //i
    .io_inputB              (pes_10_13_io_outputB[7:0]   ), //i
    .io_inputC              (pes_10_13_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_11_13), //i
    .io_outputA             (pes_11_13_io_outputA[7:0]   ), //o
    .io_outputB             (pes_11_13_io_outputB[7:0]   ), //o
    .io_outputC             (pes_11_13_io_outputC[19:0]  ), //o
    .clk                    (clk                         ), //i
    .reset                  (reset                       )  //i
  );
  ProcessingElement_144 pes_11_14 (
    .io_inputA              (pes_11_13_io_outputA[7:0]   ), //i
    .io_inputB              (pes_10_14_io_outputB[7:0]   ), //i
    .io_inputC              (pes_10_14_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_11_14), //i
    .io_outputA             (pes_11_14_io_outputA[7:0]   ), //o
    .io_outputB             (pes_11_14_io_outputB[7:0]   ), //o
    .io_outputC             (pes_11_14_io_outputC[19:0]  ), //o
    .clk                    (clk                         ), //i
    .reset                  (reset                       )  //i
  );
  ProcessingElement_159 pes_11_15 (
    .io_inputA              (pes_11_14_io_outputA[7:0]   ), //i
    .io_inputB              (pes_10_15_io_outputB[7:0]   ), //i
    .io_inputC              (pes_10_15_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_11_15), //i
    .io_outputB             (pes_11_15_io_outputB[7:0]   ), //o
    .io_outputC             (pes_11_15_io_outputC[19:0]  ), //o
    .clk                    (clk                         ), //i
    .reset                  (reset                       )  //i
  );
  ProcessingElement_144 pes_12_0 (
    .io_inputA              (skewBuffer_io_output_12[7:0]), //i
    .io_inputB              (pes_11_0_io_outputB[7:0]    ), //i
    .io_inputC              (pes_11_0_io_outputC[19:0]   ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_12_0 ), //i
    .io_outputA             (pes_12_0_io_outputA[7:0]    ), //o
    .io_outputB             (pes_12_0_io_outputB[7:0]    ), //o
    .io_outputC             (pes_12_0_io_outputC[19:0]   ), //o
    .clk                    (clk                         ), //i
    .reset                  (reset                       )  //i
  );
  ProcessingElement_144 pes_12_1 (
    .io_inputA              (pes_12_0_io_outputA[7:0]   ), //i
    .io_inputB              (pes_11_1_io_outputB[7:0]   ), //i
    .io_inputC              (pes_11_1_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_12_1), //i
    .io_outputA             (pes_12_1_io_outputA[7:0]   ), //o
    .io_outputB             (pes_12_1_io_outputB[7:0]   ), //o
    .io_outputC             (pes_12_1_io_outputC[19:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_144 pes_12_2 (
    .io_inputA              (pes_12_1_io_outputA[7:0]   ), //i
    .io_inputB              (pes_11_2_io_outputB[7:0]   ), //i
    .io_inputC              (pes_11_2_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_12_2), //i
    .io_outputA             (pes_12_2_io_outputA[7:0]   ), //o
    .io_outputB             (pes_12_2_io_outputB[7:0]   ), //o
    .io_outputC             (pes_12_2_io_outputC[19:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_144 pes_12_3 (
    .io_inputA              (pes_12_2_io_outputA[7:0]   ), //i
    .io_inputB              (pes_11_3_io_outputB[7:0]   ), //i
    .io_inputC              (pes_11_3_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_12_3), //i
    .io_outputA             (pes_12_3_io_outputA[7:0]   ), //o
    .io_outputB             (pes_12_3_io_outputB[7:0]   ), //o
    .io_outputC             (pes_12_3_io_outputC[19:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_144 pes_12_4 (
    .io_inputA              (pes_12_3_io_outputA[7:0]   ), //i
    .io_inputB              (pes_11_4_io_outputB[7:0]   ), //i
    .io_inputC              (pes_11_4_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_12_4), //i
    .io_outputA             (pes_12_4_io_outputA[7:0]   ), //o
    .io_outputB             (pes_12_4_io_outputB[7:0]   ), //o
    .io_outputC             (pes_12_4_io_outputC[19:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_144 pes_12_5 (
    .io_inputA              (pes_12_4_io_outputA[7:0]   ), //i
    .io_inputB              (pes_11_5_io_outputB[7:0]   ), //i
    .io_inputC              (pes_11_5_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_12_5), //i
    .io_outputA             (pes_12_5_io_outputA[7:0]   ), //o
    .io_outputB             (pes_12_5_io_outputB[7:0]   ), //o
    .io_outputC             (pes_12_5_io_outputC[19:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_144 pes_12_6 (
    .io_inputA              (pes_12_5_io_outputA[7:0]   ), //i
    .io_inputB              (pes_11_6_io_outputB[7:0]   ), //i
    .io_inputC              (pes_11_6_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_12_6), //i
    .io_outputA             (pes_12_6_io_outputA[7:0]   ), //o
    .io_outputB             (pes_12_6_io_outputB[7:0]   ), //o
    .io_outputC             (pes_12_6_io_outputC[19:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_144 pes_12_7 (
    .io_inputA              (pes_12_6_io_outputA[7:0]   ), //i
    .io_inputB              (pes_11_7_io_outputB[7:0]   ), //i
    .io_inputC              (pes_11_7_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_12_7), //i
    .io_outputA             (pes_12_7_io_outputA[7:0]   ), //o
    .io_outputB             (pes_12_7_io_outputB[7:0]   ), //o
    .io_outputC             (pes_12_7_io_outputC[19:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_144 pes_12_8 (
    .io_inputA              (pes_12_7_io_outputA[7:0]   ), //i
    .io_inputB              (pes_11_8_io_outputB[7:0]   ), //i
    .io_inputC              (pes_11_8_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_12_8), //i
    .io_outputA             (pes_12_8_io_outputA[7:0]   ), //o
    .io_outputB             (pes_12_8_io_outputB[7:0]   ), //o
    .io_outputC             (pes_12_8_io_outputC[19:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_144 pes_12_9 (
    .io_inputA              (pes_12_8_io_outputA[7:0]   ), //i
    .io_inputB              (pes_11_9_io_outputB[7:0]   ), //i
    .io_inputC              (pes_11_9_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_12_9), //i
    .io_outputA             (pes_12_9_io_outputA[7:0]   ), //o
    .io_outputB             (pes_12_9_io_outputB[7:0]   ), //o
    .io_outputC             (pes_12_9_io_outputC[19:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_144 pes_12_10 (
    .io_inputA              (pes_12_9_io_outputA[7:0]    ), //i
    .io_inputB              (pes_11_10_io_outputB[7:0]   ), //i
    .io_inputC              (pes_11_10_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_12_10), //i
    .io_outputA             (pes_12_10_io_outputA[7:0]   ), //o
    .io_outputB             (pes_12_10_io_outputB[7:0]   ), //o
    .io_outputC             (pes_12_10_io_outputC[19:0]  ), //o
    .clk                    (clk                         ), //i
    .reset                  (reset                       )  //i
  );
  ProcessingElement_144 pes_12_11 (
    .io_inputA              (pes_12_10_io_outputA[7:0]   ), //i
    .io_inputB              (pes_11_11_io_outputB[7:0]   ), //i
    .io_inputC              (pes_11_11_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_12_11), //i
    .io_outputA             (pes_12_11_io_outputA[7:0]   ), //o
    .io_outputB             (pes_12_11_io_outputB[7:0]   ), //o
    .io_outputC             (pes_12_11_io_outputC[19:0]  ), //o
    .clk                    (clk                         ), //i
    .reset                  (reset                       )  //i
  );
  ProcessingElement_144 pes_12_12 (
    .io_inputA              (pes_12_11_io_outputA[7:0]   ), //i
    .io_inputB              (pes_11_12_io_outputB[7:0]   ), //i
    .io_inputC              (pes_11_12_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_12_12), //i
    .io_outputA             (pes_12_12_io_outputA[7:0]   ), //o
    .io_outputB             (pes_12_12_io_outputB[7:0]   ), //o
    .io_outputC             (pes_12_12_io_outputC[19:0]  ), //o
    .clk                    (clk                         ), //i
    .reset                  (reset                       )  //i
  );
  ProcessingElement_144 pes_12_13 (
    .io_inputA              (pes_12_12_io_outputA[7:0]   ), //i
    .io_inputB              (pes_11_13_io_outputB[7:0]   ), //i
    .io_inputC              (pes_11_13_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_12_13), //i
    .io_outputA             (pes_12_13_io_outputA[7:0]   ), //o
    .io_outputB             (pes_12_13_io_outputB[7:0]   ), //o
    .io_outputC             (pes_12_13_io_outputC[19:0]  ), //o
    .clk                    (clk                         ), //i
    .reset                  (reset                       )  //i
  );
  ProcessingElement_144 pes_12_14 (
    .io_inputA              (pes_12_13_io_outputA[7:0]   ), //i
    .io_inputB              (pes_11_14_io_outputB[7:0]   ), //i
    .io_inputC              (pes_11_14_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_12_14), //i
    .io_outputA             (pes_12_14_io_outputA[7:0]   ), //o
    .io_outputB             (pes_12_14_io_outputB[7:0]   ), //o
    .io_outputC             (pes_12_14_io_outputC[19:0]  ), //o
    .clk                    (clk                         ), //i
    .reset                  (reset                       )  //i
  );
  ProcessingElement_159 pes_12_15 (
    .io_inputA              (pes_12_14_io_outputA[7:0]   ), //i
    .io_inputB              (pes_11_15_io_outputB[7:0]   ), //i
    .io_inputC              (pes_11_15_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_12_15), //i
    .io_outputB             (pes_12_15_io_outputB[7:0]   ), //o
    .io_outputC             (pes_12_15_io_outputC[19:0]  ), //o
    .clk                    (clk                         ), //i
    .reset                  (reset                       )  //i
  );
  ProcessingElement_144 pes_13_0 (
    .io_inputA              (skewBuffer_io_output_13[7:0]), //i
    .io_inputB              (pes_12_0_io_outputB[7:0]    ), //i
    .io_inputC              (pes_12_0_io_outputC[19:0]   ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_13_0 ), //i
    .io_outputA             (pes_13_0_io_outputA[7:0]    ), //o
    .io_outputB             (pes_13_0_io_outputB[7:0]    ), //o
    .io_outputC             (pes_13_0_io_outputC[19:0]   ), //o
    .clk                    (clk                         ), //i
    .reset                  (reset                       )  //i
  );
  ProcessingElement_144 pes_13_1 (
    .io_inputA              (pes_13_0_io_outputA[7:0]   ), //i
    .io_inputB              (pes_12_1_io_outputB[7:0]   ), //i
    .io_inputC              (pes_12_1_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_13_1), //i
    .io_outputA             (pes_13_1_io_outputA[7:0]   ), //o
    .io_outputB             (pes_13_1_io_outputB[7:0]   ), //o
    .io_outputC             (pes_13_1_io_outputC[19:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_144 pes_13_2 (
    .io_inputA              (pes_13_1_io_outputA[7:0]   ), //i
    .io_inputB              (pes_12_2_io_outputB[7:0]   ), //i
    .io_inputC              (pes_12_2_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_13_2), //i
    .io_outputA             (pes_13_2_io_outputA[7:0]   ), //o
    .io_outputB             (pes_13_2_io_outputB[7:0]   ), //o
    .io_outputC             (pes_13_2_io_outputC[19:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_144 pes_13_3 (
    .io_inputA              (pes_13_2_io_outputA[7:0]   ), //i
    .io_inputB              (pes_12_3_io_outputB[7:0]   ), //i
    .io_inputC              (pes_12_3_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_13_3), //i
    .io_outputA             (pes_13_3_io_outputA[7:0]   ), //o
    .io_outputB             (pes_13_3_io_outputB[7:0]   ), //o
    .io_outputC             (pes_13_3_io_outputC[19:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_144 pes_13_4 (
    .io_inputA              (pes_13_3_io_outputA[7:0]   ), //i
    .io_inputB              (pes_12_4_io_outputB[7:0]   ), //i
    .io_inputC              (pes_12_4_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_13_4), //i
    .io_outputA             (pes_13_4_io_outputA[7:0]   ), //o
    .io_outputB             (pes_13_4_io_outputB[7:0]   ), //o
    .io_outputC             (pes_13_4_io_outputC[19:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_144 pes_13_5 (
    .io_inputA              (pes_13_4_io_outputA[7:0]   ), //i
    .io_inputB              (pes_12_5_io_outputB[7:0]   ), //i
    .io_inputC              (pes_12_5_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_13_5), //i
    .io_outputA             (pes_13_5_io_outputA[7:0]   ), //o
    .io_outputB             (pes_13_5_io_outputB[7:0]   ), //o
    .io_outputC             (pes_13_5_io_outputC[19:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_144 pes_13_6 (
    .io_inputA              (pes_13_5_io_outputA[7:0]   ), //i
    .io_inputB              (pes_12_6_io_outputB[7:0]   ), //i
    .io_inputC              (pes_12_6_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_13_6), //i
    .io_outputA             (pes_13_6_io_outputA[7:0]   ), //o
    .io_outputB             (pes_13_6_io_outputB[7:0]   ), //o
    .io_outputC             (pes_13_6_io_outputC[19:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_144 pes_13_7 (
    .io_inputA              (pes_13_6_io_outputA[7:0]   ), //i
    .io_inputB              (pes_12_7_io_outputB[7:0]   ), //i
    .io_inputC              (pes_12_7_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_13_7), //i
    .io_outputA             (pes_13_7_io_outputA[7:0]   ), //o
    .io_outputB             (pes_13_7_io_outputB[7:0]   ), //o
    .io_outputC             (pes_13_7_io_outputC[19:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_144 pes_13_8 (
    .io_inputA              (pes_13_7_io_outputA[7:0]   ), //i
    .io_inputB              (pes_12_8_io_outputB[7:0]   ), //i
    .io_inputC              (pes_12_8_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_13_8), //i
    .io_outputA             (pes_13_8_io_outputA[7:0]   ), //o
    .io_outputB             (pes_13_8_io_outputB[7:0]   ), //o
    .io_outputC             (pes_13_8_io_outputC[19:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_144 pes_13_9 (
    .io_inputA              (pes_13_8_io_outputA[7:0]   ), //i
    .io_inputB              (pes_12_9_io_outputB[7:0]   ), //i
    .io_inputC              (pes_12_9_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_13_9), //i
    .io_outputA             (pes_13_9_io_outputA[7:0]   ), //o
    .io_outputB             (pes_13_9_io_outputB[7:0]   ), //o
    .io_outputC             (pes_13_9_io_outputC[19:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_144 pes_13_10 (
    .io_inputA              (pes_13_9_io_outputA[7:0]    ), //i
    .io_inputB              (pes_12_10_io_outputB[7:0]   ), //i
    .io_inputC              (pes_12_10_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_13_10), //i
    .io_outputA             (pes_13_10_io_outputA[7:0]   ), //o
    .io_outputB             (pes_13_10_io_outputB[7:0]   ), //o
    .io_outputC             (pes_13_10_io_outputC[19:0]  ), //o
    .clk                    (clk                         ), //i
    .reset                  (reset                       )  //i
  );
  ProcessingElement_144 pes_13_11 (
    .io_inputA              (pes_13_10_io_outputA[7:0]   ), //i
    .io_inputB              (pes_12_11_io_outputB[7:0]   ), //i
    .io_inputC              (pes_12_11_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_13_11), //i
    .io_outputA             (pes_13_11_io_outputA[7:0]   ), //o
    .io_outputB             (pes_13_11_io_outputB[7:0]   ), //o
    .io_outputC             (pes_13_11_io_outputC[19:0]  ), //o
    .clk                    (clk                         ), //i
    .reset                  (reset                       )  //i
  );
  ProcessingElement_144 pes_13_12 (
    .io_inputA              (pes_13_11_io_outputA[7:0]   ), //i
    .io_inputB              (pes_12_12_io_outputB[7:0]   ), //i
    .io_inputC              (pes_12_12_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_13_12), //i
    .io_outputA             (pes_13_12_io_outputA[7:0]   ), //o
    .io_outputB             (pes_13_12_io_outputB[7:0]   ), //o
    .io_outputC             (pes_13_12_io_outputC[19:0]  ), //o
    .clk                    (clk                         ), //i
    .reset                  (reset                       )  //i
  );
  ProcessingElement_144 pes_13_13 (
    .io_inputA              (pes_13_12_io_outputA[7:0]   ), //i
    .io_inputB              (pes_12_13_io_outputB[7:0]   ), //i
    .io_inputC              (pes_12_13_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_13_13), //i
    .io_outputA             (pes_13_13_io_outputA[7:0]   ), //o
    .io_outputB             (pes_13_13_io_outputB[7:0]   ), //o
    .io_outputC             (pes_13_13_io_outputC[19:0]  ), //o
    .clk                    (clk                         ), //i
    .reset                  (reset                       )  //i
  );
  ProcessingElement_144 pes_13_14 (
    .io_inputA              (pes_13_13_io_outputA[7:0]   ), //i
    .io_inputB              (pes_12_14_io_outputB[7:0]   ), //i
    .io_inputC              (pes_12_14_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_13_14), //i
    .io_outputA             (pes_13_14_io_outputA[7:0]   ), //o
    .io_outputB             (pes_13_14_io_outputB[7:0]   ), //o
    .io_outputC             (pes_13_14_io_outputC[19:0]  ), //o
    .clk                    (clk                         ), //i
    .reset                  (reset                       )  //i
  );
  ProcessingElement_159 pes_13_15 (
    .io_inputA              (pes_13_14_io_outputA[7:0]   ), //i
    .io_inputB              (pes_12_15_io_outputB[7:0]   ), //i
    .io_inputC              (pes_12_15_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_13_15), //i
    .io_outputB             (pes_13_15_io_outputB[7:0]   ), //o
    .io_outputC             (pes_13_15_io_outputC[19:0]  ), //o
    .clk                    (clk                         ), //i
    .reset                  (reset                       )  //i
  );
  ProcessingElement_144 pes_14_0 (
    .io_inputA              (skewBuffer_io_output_14[7:0]), //i
    .io_inputB              (pes_13_0_io_outputB[7:0]    ), //i
    .io_inputC              (pes_13_0_io_outputC[19:0]   ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_14_0 ), //i
    .io_outputA             (pes_14_0_io_outputA[7:0]    ), //o
    .io_outputB             (pes_14_0_io_outputB[7:0]    ), //o
    .io_outputC             (pes_14_0_io_outputC[19:0]   ), //o
    .clk                    (clk                         ), //i
    .reset                  (reset                       )  //i
  );
  ProcessingElement_144 pes_14_1 (
    .io_inputA              (pes_14_0_io_outputA[7:0]   ), //i
    .io_inputB              (pes_13_1_io_outputB[7:0]   ), //i
    .io_inputC              (pes_13_1_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_14_1), //i
    .io_outputA             (pes_14_1_io_outputA[7:0]   ), //o
    .io_outputB             (pes_14_1_io_outputB[7:0]   ), //o
    .io_outputC             (pes_14_1_io_outputC[19:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_144 pes_14_2 (
    .io_inputA              (pes_14_1_io_outputA[7:0]   ), //i
    .io_inputB              (pes_13_2_io_outputB[7:0]   ), //i
    .io_inputC              (pes_13_2_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_14_2), //i
    .io_outputA             (pes_14_2_io_outputA[7:0]   ), //o
    .io_outputB             (pes_14_2_io_outputB[7:0]   ), //o
    .io_outputC             (pes_14_2_io_outputC[19:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_144 pes_14_3 (
    .io_inputA              (pes_14_2_io_outputA[7:0]   ), //i
    .io_inputB              (pes_13_3_io_outputB[7:0]   ), //i
    .io_inputC              (pes_13_3_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_14_3), //i
    .io_outputA             (pes_14_3_io_outputA[7:0]   ), //o
    .io_outputB             (pes_14_3_io_outputB[7:0]   ), //o
    .io_outputC             (pes_14_3_io_outputC[19:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_144 pes_14_4 (
    .io_inputA              (pes_14_3_io_outputA[7:0]   ), //i
    .io_inputB              (pes_13_4_io_outputB[7:0]   ), //i
    .io_inputC              (pes_13_4_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_14_4), //i
    .io_outputA             (pes_14_4_io_outputA[7:0]   ), //o
    .io_outputB             (pes_14_4_io_outputB[7:0]   ), //o
    .io_outputC             (pes_14_4_io_outputC[19:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_144 pes_14_5 (
    .io_inputA              (pes_14_4_io_outputA[7:0]   ), //i
    .io_inputB              (pes_13_5_io_outputB[7:0]   ), //i
    .io_inputC              (pes_13_5_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_14_5), //i
    .io_outputA             (pes_14_5_io_outputA[7:0]   ), //o
    .io_outputB             (pes_14_5_io_outputB[7:0]   ), //o
    .io_outputC             (pes_14_5_io_outputC[19:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_144 pes_14_6 (
    .io_inputA              (pes_14_5_io_outputA[7:0]   ), //i
    .io_inputB              (pes_13_6_io_outputB[7:0]   ), //i
    .io_inputC              (pes_13_6_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_14_6), //i
    .io_outputA             (pes_14_6_io_outputA[7:0]   ), //o
    .io_outputB             (pes_14_6_io_outputB[7:0]   ), //o
    .io_outputC             (pes_14_6_io_outputC[19:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_144 pes_14_7 (
    .io_inputA              (pes_14_6_io_outputA[7:0]   ), //i
    .io_inputB              (pes_13_7_io_outputB[7:0]   ), //i
    .io_inputC              (pes_13_7_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_14_7), //i
    .io_outputA             (pes_14_7_io_outputA[7:0]   ), //o
    .io_outputB             (pes_14_7_io_outputB[7:0]   ), //o
    .io_outputC             (pes_14_7_io_outputC[19:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_144 pes_14_8 (
    .io_inputA              (pes_14_7_io_outputA[7:0]   ), //i
    .io_inputB              (pes_13_8_io_outputB[7:0]   ), //i
    .io_inputC              (pes_13_8_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_14_8), //i
    .io_outputA             (pes_14_8_io_outputA[7:0]   ), //o
    .io_outputB             (pes_14_8_io_outputB[7:0]   ), //o
    .io_outputC             (pes_14_8_io_outputC[19:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_144 pes_14_9 (
    .io_inputA              (pes_14_8_io_outputA[7:0]   ), //i
    .io_inputB              (pes_13_9_io_outputB[7:0]   ), //i
    .io_inputC              (pes_13_9_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_14_9), //i
    .io_outputA             (pes_14_9_io_outputA[7:0]   ), //o
    .io_outputB             (pes_14_9_io_outputB[7:0]   ), //o
    .io_outputC             (pes_14_9_io_outputC[19:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_144 pes_14_10 (
    .io_inputA              (pes_14_9_io_outputA[7:0]    ), //i
    .io_inputB              (pes_13_10_io_outputB[7:0]   ), //i
    .io_inputC              (pes_13_10_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_14_10), //i
    .io_outputA             (pes_14_10_io_outputA[7:0]   ), //o
    .io_outputB             (pes_14_10_io_outputB[7:0]   ), //o
    .io_outputC             (pes_14_10_io_outputC[19:0]  ), //o
    .clk                    (clk                         ), //i
    .reset                  (reset                       )  //i
  );
  ProcessingElement_144 pes_14_11 (
    .io_inputA              (pes_14_10_io_outputA[7:0]   ), //i
    .io_inputB              (pes_13_11_io_outputB[7:0]   ), //i
    .io_inputC              (pes_13_11_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_14_11), //i
    .io_outputA             (pes_14_11_io_outputA[7:0]   ), //o
    .io_outputB             (pes_14_11_io_outputB[7:0]   ), //o
    .io_outputC             (pes_14_11_io_outputC[19:0]  ), //o
    .clk                    (clk                         ), //i
    .reset                  (reset                       )  //i
  );
  ProcessingElement_144 pes_14_12 (
    .io_inputA              (pes_14_11_io_outputA[7:0]   ), //i
    .io_inputB              (pes_13_12_io_outputB[7:0]   ), //i
    .io_inputC              (pes_13_12_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_14_12), //i
    .io_outputA             (pes_14_12_io_outputA[7:0]   ), //o
    .io_outputB             (pes_14_12_io_outputB[7:0]   ), //o
    .io_outputC             (pes_14_12_io_outputC[19:0]  ), //o
    .clk                    (clk                         ), //i
    .reset                  (reset                       )  //i
  );
  ProcessingElement_144 pes_14_13 (
    .io_inputA              (pes_14_12_io_outputA[7:0]   ), //i
    .io_inputB              (pes_13_13_io_outputB[7:0]   ), //i
    .io_inputC              (pes_13_13_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_14_13), //i
    .io_outputA             (pes_14_13_io_outputA[7:0]   ), //o
    .io_outputB             (pes_14_13_io_outputB[7:0]   ), //o
    .io_outputC             (pes_14_13_io_outputC[19:0]  ), //o
    .clk                    (clk                         ), //i
    .reset                  (reset                       )  //i
  );
  ProcessingElement_144 pes_14_14 (
    .io_inputA              (pes_14_13_io_outputA[7:0]   ), //i
    .io_inputB              (pes_13_14_io_outputB[7:0]   ), //i
    .io_inputC              (pes_13_14_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_14_14), //i
    .io_outputA             (pes_14_14_io_outputA[7:0]   ), //o
    .io_outputB             (pes_14_14_io_outputB[7:0]   ), //o
    .io_outputC             (pes_14_14_io_outputC[19:0]  ), //o
    .clk                    (clk                         ), //i
    .reset                  (reset                       )  //i
  );
  ProcessingElement_159 pes_14_15 (
    .io_inputA              (pes_14_14_io_outputA[7:0]   ), //i
    .io_inputB              (pes_13_15_io_outputB[7:0]   ), //i
    .io_inputC              (pes_13_15_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_14_15), //i
    .io_outputB             (pes_14_15_io_outputB[7:0]   ), //o
    .io_outputC             (pes_14_15_io_outputC[19:0]  ), //o
    .clk                    (clk                         ), //i
    .reset                  (reset                       )  //i
  );
  ProcessingElement_240 pes_15_0 (
    .io_inputA              (skewBuffer_io_output_15[7:0]), //i
    .io_inputB              (pes_14_0_io_outputB[7:0]    ), //i
    .io_inputC              (pes_14_0_io_outputC[19:0]   ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_15_0 ), //i
    .io_outputA             (pes_15_0_io_outputA[7:0]    ), //o
    .io_outputC             (pes_15_0_io_outputC[19:0]   ), //o
    .clk                    (clk                         ), //i
    .reset                  (reset                       )  //i
  );
  ProcessingElement_240 pes_15_1 (
    .io_inputA              (pes_15_0_io_outputA[7:0]   ), //i
    .io_inputB              (pes_14_1_io_outputB[7:0]   ), //i
    .io_inputC              (pes_14_1_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_15_1), //i
    .io_outputA             (pes_15_1_io_outputA[7:0]   ), //o
    .io_outputC             (pes_15_1_io_outputC[19:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_240 pes_15_2 (
    .io_inputA              (pes_15_1_io_outputA[7:0]   ), //i
    .io_inputB              (pes_14_2_io_outputB[7:0]   ), //i
    .io_inputC              (pes_14_2_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_15_2), //i
    .io_outputA             (pes_15_2_io_outputA[7:0]   ), //o
    .io_outputC             (pes_15_2_io_outputC[19:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_240 pes_15_3 (
    .io_inputA              (pes_15_2_io_outputA[7:0]   ), //i
    .io_inputB              (pes_14_3_io_outputB[7:0]   ), //i
    .io_inputC              (pes_14_3_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_15_3), //i
    .io_outputA             (pes_15_3_io_outputA[7:0]   ), //o
    .io_outputC             (pes_15_3_io_outputC[19:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_240 pes_15_4 (
    .io_inputA              (pes_15_3_io_outputA[7:0]   ), //i
    .io_inputB              (pes_14_4_io_outputB[7:0]   ), //i
    .io_inputC              (pes_14_4_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_15_4), //i
    .io_outputA             (pes_15_4_io_outputA[7:0]   ), //o
    .io_outputC             (pes_15_4_io_outputC[19:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_240 pes_15_5 (
    .io_inputA              (pes_15_4_io_outputA[7:0]   ), //i
    .io_inputB              (pes_14_5_io_outputB[7:0]   ), //i
    .io_inputC              (pes_14_5_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_15_5), //i
    .io_outputA             (pes_15_5_io_outputA[7:0]   ), //o
    .io_outputC             (pes_15_5_io_outputC[19:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_240 pes_15_6 (
    .io_inputA              (pes_15_5_io_outputA[7:0]   ), //i
    .io_inputB              (pes_14_6_io_outputB[7:0]   ), //i
    .io_inputC              (pes_14_6_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_15_6), //i
    .io_outputA             (pes_15_6_io_outputA[7:0]   ), //o
    .io_outputC             (pes_15_6_io_outputC[19:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_240 pes_15_7 (
    .io_inputA              (pes_15_6_io_outputA[7:0]   ), //i
    .io_inputB              (pes_14_7_io_outputB[7:0]   ), //i
    .io_inputC              (pes_14_7_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_15_7), //i
    .io_outputA             (pes_15_7_io_outputA[7:0]   ), //o
    .io_outputC             (pes_15_7_io_outputC[19:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_240 pes_15_8 (
    .io_inputA              (pes_15_7_io_outputA[7:0]   ), //i
    .io_inputB              (pes_14_8_io_outputB[7:0]   ), //i
    .io_inputC              (pes_14_8_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_15_8), //i
    .io_outputA             (pes_15_8_io_outputA[7:0]   ), //o
    .io_outputC             (pes_15_8_io_outputC[19:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_240 pes_15_9 (
    .io_inputA              (pes_15_8_io_outputA[7:0]   ), //i
    .io_inputB              (pes_14_9_io_outputB[7:0]   ), //i
    .io_inputC              (pes_14_9_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_15_9), //i
    .io_outputA             (pes_15_9_io_outputA[7:0]   ), //o
    .io_outputC             (pes_15_9_io_outputC[19:0]  ), //o
    .clk                    (clk                        ), //i
    .reset                  (reset                      )  //i
  );
  ProcessingElement_240 pes_15_10 (
    .io_inputA              (pes_15_9_io_outputA[7:0]    ), //i
    .io_inputB              (pes_14_10_io_outputB[7:0]   ), //i
    .io_inputC              (pes_14_10_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_15_10), //i
    .io_outputA             (pes_15_10_io_outputA[7:0]   ), //o
    .io_outputC             (pes_15_10_io_outputC[19:0]  ), //o
    .clk                    (clk                         ), //i
    .reset                  (reset                       )  //i
  );
  ProcessingElement_240 pes_15_11 (
    .io_inputA              (pes_15_10_io_outputA[7:0]   ), //i
    .io_inputB              (pes_14_11_io_outputB[7:0]   ), //i
    .io_inputC              (pes_14_11_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_15_11), //i
    .io_outputA             (pes_15_11_io_outputA[7:0]   ), //o
    .io_outputC             (pes_15_11_io_outputC[19:0]  ), //o
    .clk                    (clk                         ), //i
    .reset                  (reset                       )  //i
  );
  ProcessingElement_240 pes_15_12 (
    .io_inputA              (pes_15_11_io_outputA[7:0]   ), //i
    .io_inputB              (pes_14_12_io_outputB[7:0]   ), //i
    .io_inputC              (pes_14_12_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_15_12), //i
    .io_outputA             (pes_15_12_io_outputA[7:0]   ), //o
    .io_outputC             (pes_15_12_io_outputC[19:0]  ), //o
    .clk                    (clk                         ), //i
    .reset                  (reset                       )  //i
  );
  ProcessingElement_240 pes_15_13 (
    .io_inputA              (pes_15_12_io_outputA[7:0]   ), //i
    .io_inputB              (pes_14_13_io_outputB[7:0]   ), //i
    .io_inputC              (pes_14_13_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_15_13), //i
    .io_outputA             (pes_15_13_io_outputA[7:0]   ), //o
    .io_outputC             (pes_15_13_io_outputC[19:0]  ), //o
    .clk                    (clk                         ), //i
    .reset                  (reset                       )  //i
  );
  ProcessingElement_240 pes_15_14 (
    .io_inputA              (pes_15_13_io_outputA[7:0]   ), //i
    .io_inputB              (pes_14_14_io_outputB[7:0]   ), //i
    .io_inputC              (pes_14_14_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_15_14), //i
    .io_outputA             (pes_15_14_io_outputA[7:0]   ), //o
    .io_outputC             (pes_15_14_io_outputC[19:0]  ), //o
    .clk                    (clk                         ), //i
    .reset                  (reset                       )  //i
  );
  ProcessingElement_255 pes_15_15 (
    .io_inputA              (pes_15_14_io_outputA[7:0]   ), //i
    .io_inputB              (pes_14_15_io_outputB[7:0]   ), //i
    .io_inputC              (pes_14_15_io_outputC[19:0]  ), //i
    .io_inputCaptureEnableB (io_inputCaptureEnableB_15_15), //i
    .io_outputC             (pes_15_15_io_outputC[19:0]  ), //o
    .clk                    (clk                         ), //i
    .reset                  (reset                       )  //i
  );
//#endregion

//#region Skew Buffer
  TypeA_SkewBuffer skewBuffer (
    .io_input_0   (io_inputA_0[7:0]            ), //i
    .io_input_1   (io_inputA_1[7:0]            ), //i
    .io_input_2   (io_inputA_2[7:0]            ), //i
    .io_input_3   (io_inputA_3[7:0]            ), //i
    .io_input_4   (io_inputA_4[7:0]            ), //i
    .io_input_5   (io_inputA_5[7:0]            ), //i
    .io_input_6   (io_inputA_6[7:0]            ), //i
    .io_input_7   (io_inputA_7[7:0]            ), //i
    .io_input_8   (io_inputA_8[7:0]            ), //i
    .io_input_9   (io_inputA_9[7:0]            ), //i
    .io_input_10  (io_inputA_10[7:0]           ), //i
    .io_input_11  (io_inputA_11[7:0]           ), //i
    .io_input_12  (io_inputA_12[7:0]           ), //i
    .io_input_13  (io_inputA_13[7:0]           ), //i
    .io_input_14  (io_inputA_14[7:0]           ), //i
    .io_input_15  (io_inputA_15[7:0]           ), //i
    .io_output_0  (skewBuffer_io_output_0[7:0] ), //o
    .io_output_1  (skewBuffer_io_output_1[7:0] ), //o
    .io_output_2  (skewBuffer_io_output_2[7:0] ), //o
    .io_output_3  (skewBuffer_io_output_3[7:0] ), //o
    .io_output_4  (skewBuffer_io_output_4[7:0] ), //o
    .io_output_5  (skewBuffer_io_output_5[7:0] ), //o
    .io_output_6  (skewBuffer_io_output_6[7:0] ), //o
    .io_output_7  (skewBuffer_io_output_7[7:0] ), //o
    .io_output_8  (skewBuffer_io_output_8[7:0] ), //o
    .io_output_9  (skewBuffer_io_output_9[7:0] ), //o
    .io_output_10 (skewBuffer_io_output_10[7:0]), //o
    .io_output_11 (skewBuffer_io_output_11[7:0]), //o
    .io_output_12 (skewBuffer_io_output_12[7:0]), //o
    .io_output_13 (skewBuffer_io_output_13[7:0]), //o
    .io_output_14 (skewBuffer_io_output_14[7:0]), //o
    .io_output_15 (skewBuffer_io_output_15[7:0]), //o
    .clk          (clk                         ), //i
    .reset        (reset                       )  //i
  );
  TypeC_DeskewBuffer skewBuffer_1 (
    .io_input_0   (pes_15_0_io_outputC[19:0]      ), //i
    .io_input_1   (pes_15_1_io_outputC[19:0]      ), //i
    .io_input_2   (pes_15_2_io_outputC[19:0]      ), //i
    .io_input_3   (pes_15_3_io_outputC[19:0]      ), //i
    .io_input_4   (pes_15_4_io_outputC[19:0]      ), //i
    .io_input_5   (pes_15_5_io_outputC[19:0]      ), //i
    .io_input_6   (pes_15_6_io_outputC[19:0]      ), //i
    .io_input_7   (pes_15_7_io_outputC[19:0]      ), //i
    .io_input_8   (pes_15_8_io_outputC[19:0]      ), //i
    .io_input_9   (pes_15_9_io_outputC[19:0]      ), //i
    .io_input_10  (pes_15_10_io_outputC[19:0]     ), //i
    .io_input_11  (pes_15_11_io_outputC[19:0]     ), //i
    .io_input_12  (pes_15_12_io_outputC[19:0]     ), //i
    .io_input_13  (pes_15_13_io_outputC[19:0]     ), //i
    .io_input_14  (pes_15_14_io_outputC[19:0]     ), //i
    .io_input_15  (pes_15_15_io_outputC[19:0]     ), //i
    .io_output_0  (skewBuffer_1_io_output_0[19:0] ), //o
    .io_output_1  (skewBuffer_1_io_output_1[19:0] ), //o
    .io_output_2  (skewBuffer_1_io_output_2[19:0] ), //o
    .io_output_3  (skewBuffer_1_io_output_3[19:0] ), //o
    .io_output_4  (skewBuffer_1_io_output_4[19:0] ), //o
    .io_output_5  (skewBuffer_1_io_output_5[19:0] ), //o
    .io_output_6  (skewBuffer_1_io_output_6[19:0] ), //o
    .io_output_7  (skewBuffer_1_io_output_7[19:0] ), //o
    .io_output_8  (skewBuffer_1_io_output_8[19:0] ), //o
    .io_output_9  (skewBuffer_1_io_output_9[19:0] ), //o
    .io_output_10 (skewBuffer_1_io_output_10[19:0]), //o
    .io_output_11 (skewBuffer_1_io_output_11[19:0]), //o
    .io_output_12 (skewBuffer_1_io_output_12[19:0]), //o
    .io_output_13 (skewBuffer_1_io_output_13[19:0]), //o
    .io_output_14 (skewBuffer_1_io_output_14[19:0]), //o
    .io_output_15 (skewBuffer_1_io_output_15[19:0]), //o
    .clk          (clk                            ), //i
    .reset        (reset                          )  //i
  );
//#endregion

//#region Assignments
  assign io_outputC_0 = skewBuffer_1_io_output_0;
  assign io_outputC_1 = skewBuffer_1_io_output_1;
  assign io_outputC_2 = skewBuffer_1_io_output_2;
  assign io_outputC_3 = skewBuffer_1_io_output_3;
  assign io_outputC_4 = skewBuffer_1_io_output_4;
  assign io_outputC_5 = skewBuffer_1_io_output_5;
  assign io_outputC_6 = skewBuffer_1_io_output_6;
  assign io_outputC_7 = skewBuffer_1_io_output_7;
  assign io_outputC_8 = skewBuffer_1_io_output_8;
  assign io_outputC_9 = skewBuffer_1_io_output_9;
  assign io_outputC_10 = skewBuffer_1_io_output_10;
  assign io_outputC_11 = skewBuffer_1_io_output_11;
  assign io_outputC_12 = skewBuffer_1_io_output_12;
  assign io_outputC_13 = skewBuffer_1_io_output_13;
  assign io_outputC_14 = skewBuffer_1_io_output_14;
  assign io_outputC_15 = skewBuffer_1_io_output_15;
  always @(posedge clk) begin
    io_inputB_0_regNext <= io_inputB_0;
    io_inputB_1_regNext <= io_inputB_1;
    io_inputB_2_regNext <= io_inputB_2;
    io_inputB_3_regNext <= io_inputB_3;
    io_inputB_4_regNext <= io_inputB_4;
    io_inputB_5_regNext <= io_inputB_5;
    io_inputB_6_regNext <= io_inputB_6;
    io_inputB_7_regNext <= io_inputB_7;
    io_inputB_8_regNext <= io_inputB_8;
    io_inputB_9_regNext <= io_inputB_9;
    io_inputB_10_regNext <= io_inputB_10;
    io_inputB_11_regNext <= io_inputB_11;
    io_inputB_12_regNext <= io_inputB_12;
    io_inputB_13_regNext <= io_inputB_13;
    io_inputB_14_regNext <= io_inputB_14;
    io_inputB_15_regNext <= io_inputB_15;
  end
//#endregion

endmodule

module TypeC_DeskewBuffer (
  input  wire [19:0]   io_input_0,
  input  wire [19:0]   io_input_1,
  input  wire [19:0]   io_input_2,
  input  wire [19:0]   io_input_3,
  input  wire [19:0]   io_input_4,
  input  wire [19:0]   io_input_5,
  input  wire [19:0]   io_input_6,
  input  wire [19:0]   io_input_7,
  input  wire [19:0]   io_input_8,
  input  wire [19:0]   io_input_9,
  input  wire [19:0]   io_input_10,
  input  wire [19:0]   io_input_11,
  input  wire [19:0]   io_input_12,
  input  wire [19:0]   io_input_13,
  input  wire [19:0]   io_input_14,
  input  wire [19:0]   io_input_15,
  output wire [19:0]   io_output_0,
  output wire [19:0]   io_output_1,
  output wire [19:0]   io_output_2,
  output wire [19:0]   io_output_3,
  output wire [19:0]   io_output_4,
  output wire [19:0]   io_output_5,
  output wire [19:0]   io_output_6,
  output wire [19:0]   io_output_7,
  output wire [19:0]   io_output_8,
  output wire [19:0]   io_output_9,
  output wire [19:0]   io_output_10,
  output wire [19:0]   io_output_11,
  output wire [19:0]   io_output_12,
  output wire [19:0]   io_output_13,
  output wire [19:0]   io_output_14,
  output wire [19:0]   io_output_15,
  input  wire          clk,
  input  wire          reset
);

  reg        [19:0]   io_input_0_delay_1;
  reg        [19:0]   io_input_0_delay_2;
  reg        [19:0]   io_input_0_delay_3;
  reg        [19:0]   io_input_0_delay_4;
  reg        [19:0]   io_input_0_delay_5;
  reg        [19:0]   io_input_0_delay_6;
  reg        [19:0]   io_input_0_delay_7;
  reg        [19:0]   io_input_0_delay_8;
  reg        [19:0]   io_input_0_delay_9;
  reg        [19:0]   io_input_0_delay_10;
  reg        [19:0]   io_input_0_delay_11;
  reg        [19:0]   io_input_0_delay_12;
  reg        [19:0]   io_input_0_delay_13;
  reg        [19:0]   io_input_0_delay_14;
  reg        [19:0]   io_input_0_delay_15;
  reg        [19:0]   io_input_0_delay_16;
  reg        [19:0]   io_input_1_delay_1;
  reg        [19:0]   io_input_1_delay_2;
  reg        [19:0]   io_input_1_delay_3;
  reg        [19:0]   io_input_1_delay_4;
  reg        [19:0]   io_input_1_delay_5;
  reg        [19:0]   io_input_1_delay_6;
  reg        [19:0]   io_input_1_delay_7;
  reg        [19:0]   io_input_1_delay_8;
  reg        [19:0]   io_input_1_delay_9;
  reg        [19:0]   io_input_1_delay_10;
  reg        [19:0]   io_input_1_delay_11;
  reg        [19:0]   io_input_1_delay_12;
  reg        [19:0]   io_input_1_delay_13;
  reg        [19:0]   io_input_1_delay_14;
  reg        [19:0]   io_input_1_delay_15;
  reg        [19:0]   io_input_2_delay_1;
  reg        [19:0]   io_input_2_delay_2;
  reg        [19:0]   io_input_2_delay_3;
  reg        [19:0]   io_input_2_delay_4;
  reg        [19:0]   io_input_2_delay_5;
  reg        [19:0]   io_input_2_delay_6;
  reg        [19:0]   io_input_2_delay_7;
  reg        [19:0]   io_input_2_delay_8;
  reg        [19:0]   io_input_2_delay_9;
  reg        [19:0]   io_input_2_delay_10;
  reg        [19:0]   io_input_2_delay_11;
  reg        [19:0]   io_input_2_delay_12;
  reg        [19:0]   io_input_2_delay_13;
  reg        [19:0]   io_input_2_delay_14;
  reg        [19:0]   io_input_3_delay_1;
  reg        [19:0]   io_input_3_delay_2;
  reg        [19:0]   io_input_3_delay_3;
  reg        [19:0]   io_input_3_delay_4;
  reg        [19:0]   io_input_3_delay_5;
  reg        [19:0]   io_input_3_delay_6;
  reg        [19:0]   io_input_3_delay_7;
  reg        [19:0]   io_input_3_delay_8;
  reg        [19:0]   io_input_3_delay_9;
  reg        [19:0]   io_input_3_delay_10;
  reg        [19:0]   io_input_3_delay_11;
  reg        [19:0]   io_input_3_delay_12;
  reg        [19:0]   io_input_3_delay_13;
  reg        [19:0]   io_input_4_delay_1;
  reg        [19:0]   io_input_4_delay_2;
  reg        [19:0]   io_input_4_delay_3;
  reg        [19:0]   io_input_4_delay_4;
  reg        [19:0]   io_input_4_delay_5;
  reg        [19:0]   io_input_4_delay_6;
  reg        [19:0]   io_input_4_delay_7;
  reg        [19:0]   io_input_4_delay_8;
  reg        [19:0]   io_input_4_delay_9;
  reg        [19:0]   io_input_4_delay_10;
  reg        [19:0]   io_input_4_delay_11;
  reg        [19:0]   io_input_4_delay_12;
  reg        [19:0]   io_input_5_delay_1;
  reg        [19:0]   io_input_5_delay_2;
  reg        [19:0]   io_input_5_delay_3;
  reg        [19:0]   io_input_5_delay_4;
  reg        [19:0]   io_input_5_delay_5;
  reg        [19:0]   io_input_5_delay_6;
  reg        [19:0]   io_input_5_delay_7;
  reg        [19:0]   io_input_5_delay_8;
  reg        [19:0]   io_input_5_delay_9;
  reg        [19:0]   io_input_5_delay_10;
  reg        [19:0]   io_input_5_delay_11;
  reg        [19:0]   io_input_6_delay_1;
  reg        [19:0]   io_input_6_delay_2;
  reg        [19:0]   io_input_6_delay_3;
  reg        [19:0]   io_input_6_delay_4;
  reg        [19:0]   io_input_6_delay_5;
  reg        [19:0]   io_input_6_delay_6;
  reg        [19:0]   io_input_6_delay_7;
  reg        [19:0]   io_input_6_delay_8;
  reg        [19:0]   io_input_6_delay_9;
  reg        [19:0]   io_input_6_delay_10;
  reg        [19:0]   io_input_7_delay_1;
  reg        [19:0]   io_input_7_delay_2;
  reg        [19:0]   io_input_7_delay_3;
  reg        [19:0]   io_input_7_delay_4;
  reg        [19:0]   io_input_7_delay_5;
  reg        [19:0]   io_input_7_delay_6;
  reg        [19:0]   io_input_7_delay_7;
  reg        [19:0]   io_input_7_delay_8;
  reg        [19:0]   io_input_7_delay_9;
  reg        [19:0]   io_input_8_delay_1;
  reg        [19:0]   io_input_8_delay_2;
  reg        [19:0]   io_input_8_delay_3;
  reg        [19:0]   io_input_8_delay_4;
  reg        [19:0]   io_input_8_delay_5;
  reg        [19:0]   io_input_8_delay_6;
  reg        [19:0]   io_input_8_delay_7;
  reg        [19:0]   io_input_8_delay_8;
  reg        [19:0]   io_input_9_delay_1;
  reg        [19:0]   io_input_9_delay_2;
  reg        [19:0]   io_input_9_delay_3;
  reg        [19:0]   io_input_9_delay_4;
  reg        [19:0]   io_input_9_delay_5;
  reg        [19:0]   io_input_9_delay_6;
  reg        [19:0]   io_input_9_delay_7;
  reg        [19:0]   io_input_10_delay_1;
  reg        [19:0]   io_input_10_delay_2;
  reg        [19:0]   io_input_10_delay_3;
  reg        [19:0]   io_input_10_delay_4;
  reg        [19:0]   io_input_10_delay_5;
  reg        [19:0]   io_input_10_delay_6;
  reg        [19:0]   io_input_11_delay_1;
  reg        [19:0]   io_input_11_delay_2;
  reg        [19:0]   io_input_11_delay_3;
  reg        [19:0]   io_input_11_delay_4;
  reg        [19:0]   io_input_11_delay_5;
  reg        [19:0]   io_input_12_delay_1;
  reg        [19:0]   io_input_12_delay_2;
  reg        [19:0]   io_input_12_delay_3;
  reg        [19:0]   io_input_12_delay_4;
  reg        [19:0]   io_input_13_delay_1;
  reg        [19:0]   io_input_13_delay_2;
  reg        [19:0]   io_input_13_delay_3;
  reg        [19:0]   io_input_14_delay_1;
  reg        [19:0]   io_input_14_delay_2;
  reg        [19:0]   io_input_15_delay_1;

  assign io_output_0 = io_input_0_delay_16;
  assign io_output_1 = io_input_1_delay_15;
  assign io_output_2 = io_input_2_delay_14;
  assign io_output_3 = io_input_3_delay_13;
  assign io_output_4 = io_input_4_delay_12;
  assign io_output_5 = io_input_5_delay_11;
  assign io_output_6 = io_input_6_delay_10;
  assign io_output_7 = io_input_7_delay_9;
  assign io_output_8 = io_input_8_delay_8;
  assign io_output_9 = io_input_9_delay_7;
  assign io_output_10 = io_input_10_delay_6;
  assign io_output_11 = io_input_11_delay_5;
  assign io_output_12 = io_input_12_delay_4;
  assign io_output_13 = io_input_13_delay_3;
  assign io_output_14 = io_input_14_delay_2;
  assign io_output_15 = io_input_15_delay_1;
  always @(posedge clk) begin
    io_input_0_delay_1 <= io_input_0;
    io_input_0_delay_2 <= io_input_0_delay_1;
    io_input_0_delay_3 <= io_input_0_delay_2;
    io_input_0_delay_4 <= io_input_0_delay_3;
    io_input_0_delay_5 <= io_input_0_delay_4;
    io_input_0_delay_6 <= io_input_0_delay_5;
    io_input_0_delay_7 <= io_input_0_delay_6;
    io_input_0_delay_8 <= io_input_0_delay_7;
    io_input_0_delay_9 <= io_input_0_delay_8;
    io_input_0_delay_10 <= io_input_0_delay_9;
    io_input_0_delay_11 <= io_input_0_delay_10;
    io_input_0_delay_12 <= io_input_0_delay_11;
    io_input_0_delay_13 <= io_input_0_delay_12;
    io_input_0_delay_14 <= io_input_0_delay_13;
    io_input_0_delay_15 <= io_input_0_delay_14;
    io_input_0_delay_16 <= io_input_0_delay_15;
    io_input_1_delay_1 <= io_input_1;
    io_input_1_delay_2 <= io_input_1_delay_1;
    io_input_1_delay_3 <= io_input_1_delay_2;
    io_input_1_delay_4 <= io_input_1_delay_3;
    io_input_1_delay_5 <= io_input_1_delay_4;
    io_input_1_delay_6 <= io_input_1_delay_5;
    io_input_1_delay_7 <= io_input_1_delay_6;
    io_input_1_delay_8 <= io_input_1_delay_7;
    io_input_1_delay_9 <= io_input_1_delay_8;
    io_input_1_delay_10 <= io_input_1_delay_9;
    io_input_1_delay_11 <= io_input_1_delay_10;
    io_input_1_delay_12 <= io_input_1_delay_11;
    io_input_1_delay_13 <= io_input_1_delay_12;
    io_input_1_delay_14 <= io_input_1_delay_13;
    io_input_1_delay_15 <= io_input_1_delay_14;
    io_input_2_delay_1 <= io_input_2;
    io_input_2_delay_2 <= io_input_2_delay_1;
    io_input_2_delay_3 <= io_input_2_delay_2;
    io_input_2_delay_4 <= io_input_2_delay_3;
    io_input_2_delay_5 <= io_input_2_delay_4;
    io_input_2_delay_6 <= io_input_2_delay_5;
    io_input_2_delay_7 <= io_input_2_delay_6;
    io_input_2_delay_8 <= io_input_2_delay_7;
    io_input_2_delay_9 <= io_input_2_delay_8;
    io_input_2_delay_10 <= io_input_2_delay_9;
    io_input_2_delay_11 <= io_input_2_delay_10;
    io_input_2_delay_12 <= io_input_2_delay_11;
    io_input_2_delay_13 <= io_input_2_delay_12;
    io_input_2_delay_14 <= io_input_2_delay_13;
    io_input_3_delay_1 <= io_input_3;
    io_input_3_delay_2 <= io_input_3_delay_1;
    io_input_3_delay_3 <= io_input_3_delay_2;
    io_input_3_delay_4 <= io_input_3_delay_3;
    io_input_3_delay_5 <= io_input_3_delay_4;
    io_input_3_delay_6 <= io_input_3_delay_5;
    io_input_3_delay_7 <= io_input_3_delay_6;
    io_input_3_delay_8 <= io_input_3_delay_7;
    io_input_3_delay_9 <= io_input_3_delay_8;
    io_input_3_delay_10 <= io_input_3_delay_9;
    io_input_3_delay_11 <= io_input_3_delay_10;
    io_input_3_delay_12 <= io_input_3_delay_11;
    io_input_3_delay_13 <= io_input_3_delay_12;
    io_input_4_delay_1 <= io_input_4;
    io_input_4_delay_2 <= io_input_4_delay_1;
    io_input_4_delay_3 <= io_input_4_delay_2;
    io_input_4_delay_4 <= io_input_4_delay_3;
    io_input_4_delay_5 <= io_input_4_delay_4;
    io_input_4_delay_6 <= io_input_4_delay_5;
    io_input_4_delay_7 <= io_input_4_delay_6;
    io_input_4_delay_8 <= io_input_4_delay_7;
    io_input_4_delay_9 <= io_input_4_delay_8;
    io_input_4_delay_10 <= io_input_4_delay_9;
    io_input_4_delay_11 <= io_input_4_delay_10;
    io_input_4_delay_12 <= io_input_4_delay_11;
    io_input_5_delay_1 <= io_input_5;
    io_input_5_delay_2 <= io_input_5_delay_1;
    io_input_5_delay_3 <= io_input_5_delay_2;
    io_input_5_delay_4 <= io_input_5_delay_3;
    io_input_5_delay_5 <= io_input_5_delay_4;
    io_input_5_delay_6 <= io_input_5_delay_5;
    io_input_5_delay_7 <= io_input_5_delay_6;
    io_input_5_delay_8 <= io_input_5_delay_7;
    io_input_5_delay_9 <= io_input_5_delay_8;
    io_input_5_delay_10 <= io_input_5_delay_9;
    io_input_5_delay_11 <= io_input_5_delay_10;
    io_input_6_delay_1 <= io_input_6;
    io_input_6_delay_2 <= io_input_6_delay_1;
    io_input_6_delay_3 <= io_input_6_delay_2;
    io_input_6_delay_4 <= io_input_6_delay_3;
    io_input_6_delay_5 <= io_input_6_delay_4;
    io_input_6_delay_6 <= io_input_6_delay_5;
    io_input_6_delay_7 <= io_input_6_delay_6;
    io_input_6_delay_8 <= io_input_6_delay_7;
    io_input_6_delay_9 <= io_input_6_delay_8;
    io_input_6_delay_10 <= io_input_6_delay_9;
    io_input_7_delay_1 <= io_input_7;
    io_input_7_delay_2 <= io_input_7_delay_1;
    io_input_7_delay_3 <= io_input_7_delay_2;
    io_input_7_delay_4 <= io_input_7_delay_3;
    io_input_7_delay_5 <= io_input_7_delay_4;
    io_input_7_delay_6 <= io_input_7_delay_5;
    io_input_7_delay_7 <= io_input_7_delay_6;
    io_input_7_delay_8 <= io_input_7_delay_7;
    io_input_7_delay_9 <= io_input_7_delay_8;
    io_input_8_delay_1 <= io_input_8;
    io_input_8_delay_2 <= io_input_8_delay_1;
    io_input_8_delay_3 <= io_input_8_delay_2;
    io_input_8_delay_4 <= io_input_8_delay_3;
    io_input_8_delay_5 <= io_input_8_delay_4;
    io_input_8_delay_6 <= io_input_8_delay_5;
    io_input_8_delay_7 <= io_input_8_delay_6;
    io_input_8_delay_8 <= io_input_8_delay_7;
    io_input_9_delay_1 <= io_input_9;
    io_input_9_delay_2 <= io_input_9_delay_1;
    io_input_9_delay_3 <= io_input_9_delay_2;
    io_input_9_delay_4 <= io_input_9_delay_3;
    io_input_9_delay_5 <= io_input_9_delay_4;
    io_input_9_delay_6 <= io_input_9_delay_5;
    io_input_9_delay_7 <= io_input_9_delay_6;
    io_input_10_delay_1 <= io_input_10;
    io_input_10_delay_2 <= io_input_10_delay_1;
    io_input_10_delay_3 <= io_input_10_delay_2;
    io_input_10_delay_4 <= io_input_10_delay_3;
    io_input_10_delay_5 <= io_input_10_delay_4;
    io_input_10_delay_6 <= io_input_10_delay_5;
    io_input_11_delay_1 <= io_input_11;
    io_input_11_delay_2 <= io_input_11_delay_1;
    io_input_11_delay_3 <= io_input_11_delay_2;
    io_input_11_delay_4 <= io_input_11_delay_3;
    io_input_11_delay_5 <= io_input_11_delay_4;
    io_input_12_delay_1 <= io_input_12;
    io_input_12_delay_2 <= io_input_12_delay_1;
    io_input_12_delay_3 <= io_input_12_delay_2;
    io_input_12_delay_4 <= io_input_12_delay_3;
    io_input_13_delay_1 <= io_input_13;
    io_input_13_delay_2 <= io_input_13_delay_1;
    io_input_13_delay_3 <= io_input_13_delay_2;
    io_input_14_delay_1 <= io_input_14;
    io_input_14_delay_2 <= io_input_14_delay_1;
    io_input_15_delay_1 <= io_input_15;
  end


endmodule

module TypeA_SkewBuffer (
  input  wire [7:0]    io_input_0,
  input  wire [7:0]    io_input_1,
  input  wire [7:0]    io_input_2,
  input  wire [7:0]    io_input_3,
  input  wire [7:0]    io_input_4,
  input  wire [7:0]    io_input_5,
  input  wire [7:0]    io_input_6,
  input  wire [7:0]    io_input_7,
  input  wire [7:0]    io_input_8,
  input  wire [7:0]    io_input_9,
  input  wire [7:0]    io_input_10,
  input  wire [7:0]    io_input_11,
  input  wire [7:0]    io_input_12,
  input  wire [7:0]    io_input_13,
  input  wire [7:0]    io_input_14,
  input  wire [7:0]    io_input_15,
  output wire [7:0]    io_output_0,
  output wire [7:0]    io_output_1,
  output wire [7:0]    io_output_2,
  output wire [7:0]    io_output_3,
  output wire [7:0]    io_output_4,
  output wire [7:0]    io_output_5,
  output wire [7:0]    io_output_6,
  output wire [7:0]    io_output_7,
  output wire [7:0]    io_output_8,
  output wire [7:0]    io_output_9,
  output wire [7:0]    io_output_10,
  output wire [7:0]    io_output_11,
  output wire [7:0]    io_output_12,
  output wire [7:0]    io_output_13,
  output wire [7:0]    io_output_14,
  output wire [7:0]    io_output_15,
  input  wire          clk,
  input  wire          reset
);

  reg        [7:0]    io_input_0_delay_1;
  reg        [7:0]    io_input_1_delay_1;
  reg        [7:0]    io_input_1_delay_2;
  reg        [7:0]    io_input_2_delay_1;
  reg        [7:0]    io_input_2_delay_2;
  reg        [7:0]    io_input_2_delay_3;
  reg        [7:0]    io_input_3_delay_1;
  reg        [7:0]    io_input_3_delay_2;
  reg        [7:0]    io_input_3_delay_3;
  reg        [7:0]    io_input_3_delay_4;
  reg        [7:0]    io_input_4_delay_1;
  reg        [7:0]    io_input_4_delay_2;
  reg        [7:0]    io_input_4_delay_3;
  reg        [7:0]    io_input_4_delay_4;
  reg        [7:0]    io_input_4_delay_5;
  reg        [7:0]    io_input_5_delay_1;
  reg        [7:0]    io_input_5_delay_2;
  reg        [7:0]    io_input_5_delay_3;
  reg        [7:0]    io_input_5_delay_4;
  reg        [7:0]    io_input_5_delay_5;
  reg        [7:0]    io_input_5_delay_6;
  reg        [7:0]    io_input_6_delay_1;
  reg        [7:0]    io_input_6_delay_2;
  reg        [7:0]    io_input_6_delay_3;
  reg        [7:0]    io_input_6_delay_4;
  reg        [7:0]    io_input_6_delay_5;
  reg        [7:0]    io_input_6_delay_6;
  reg        [7:0]    io_input_6_delay_7;
  reg        [7:0]    io_input_7_delay_1;
  reg        [7:0]    io_input_7_delay_2;
  reg        [7:0]    io_input_7_delay_3;
  reg        [7:0]    io_input_7_delay_4;
  reg        [7:0]    io_input_7_delay_5;
  reg        [7:0]    io_input_7_delay_6;
  reg        [7:0]    io_input_7_delay_7;
  reg        [7:0]    io_input_7_delay_8;
  reg        [7:0]    io_input_8_delay_1;
  reg        [7:0]    io_input_8_delay_2;
  reg        [7:0]    io_input_8_delay_3;
  reg        [7:0]    io_input_8_delay_4;
  reg        [7:0]    io_input_8_delay_5;
  reg        [7:0]    io_input_8_delay_6;
  reg        [7:0]    io_input_8_delay_7;
  reg        [7:0]    io_input_8_delay_8;
  reg        [7:0]    io_input_8_delay_9;
  reg        [7:0]    io_input_9_delay_1;
  reg        [7:0]    io_input_9_delay_2;
  reg        [7:0]    io_input_9_delay_3;
  reg        [7:0]    io_input_9_delay_4;
  reg        [7:0]    io_input_9_delay_5;
  reg        [7:0]    io_input_9_delay_6;
  reg        [7:0]    io_input_9_delay_7;
  reg        [7:0]    io_input_9_delay_8;
  reg        [7:0]    io_input_9_delay_9;
  reg        [7:0]    io_input_9_delay_10;
  reg        [7:0]    io_input_10_delay_1;
  reg        [7:0]    io_input_10_delay_2;
  reg        [7:0]    io_input_10_delay_3;
  reg        [7:0]    io_input_10_delay_4;
  reg        [7:0]    io_input_10_delay_5;
  reg        [7:0]    io_input_10_delay_6;
  reg        [7:0]    io_input_10_delay_7;
  reg        [7:0]    io_input_10_delay_8;
  reg        [7:0]    io_input_10_delay_9;
  reg        [7:0]    io_input_10_delay_10;
  reg        [7:0]    io_input_10_delay_11;
  reg        [7:0]    io_input_11_delay_1;
  reg        [7:0]    io_input_11_delay_2;
  reg        [7:0]    io_input_11_delay_3;
  reg        [7:0]    io_input_11_delay_4;
  reg        [7:0]    io_input_11_delay_5;
  reg        [7:0]    io_input_11_delay_6;
  reg        [7:0]    io_input_11_delay_7;
  reg        [7:0]    io_input_11_delay_8;
  reg        [7:0]    io_input_11_delay_9;
  reg        [7:0]    io_input_11_delay_10;
  reg        [7:0]    io_input_11_delay_11;
  reg        [7:0]    io_input_11_delay_12;
  reg        [7:0]    io_input_12_delay_1;
  reg        [7:0]    io_input_12_delay_2;
  reg        [7:0]    io_input_12_delay_3;
  reg        [7:0]    io_input_12_delay_4;
  reg        [7:0]    io_input_12_delay_5;
  reg        [7:0]    io_input_12_delay_6;
  reg        [7:0]    io_input_12_delay_7;
  reg        [7:0]    io_input_12_delay_8;
  reg        [7:0]    io_input_12_delay_9;
  reg        [7:0]    io_input_12_delay_10;
  reg        [7:0]    io_input_12_delay_11;
  reg        [7:0]    io_input_12_delay_12;
  reg        [7:0]    io_input_12_delay_13;
  reg        [7:0]    io_input_13_delay_1;
  reg        [7:0]    io_input_13_delay_2;
  reg        [7:0]    io_input_13_delay_3;
  reg        [7:0]    io_input_13_delay_4;
  reg        [7:0]    io_input_13_delay_5;
  reg        [7:0]    io_input_13_delay_6;
  reg        [7:0]    io_input_13_delay_7;
  reg        [7:0]    io_input_13_delay_8;
  reg        [7:0]    io_input_13_delay_9;
  reg        [7:0]    io_input_13_delay_10;
  reg        [7:0]    io_input_13_delay_11;
  reg        [7:0]    io_input_13_delay_12;
  reg        [7:0]    io_input_13_delay_13;
  reg        [7:0]    io_input_13_delay_14;
  reg        [7:0]    io_input_14_delay_1;
  reg        [7:0]    io_input_14_delay_2;
  reg        [7:0]    io_input_14_delay_3;
  reg        [7:0]    io_input_14_delay_4;
  reg        [7:0]    io_input_14_delay_5;
  reg        [7:0]    io_input_14_delay_6;
  reg        [7:0]    io_input_14_delay_7;
  reg        [7:0]    io_input_14_delay_8;
  reg        [7:0]    io_input_14_delay_9;
  reg        [7:0]    io_input_14_delay_10;
  reg        [7:0]    io_input_14_delay_11;
  reg        [7:0]    io_input_14_delay_12;
  reg        [7:0]    io_input_14_delay_13;
  reg        [7:0]    io_input_14_delay_14;
  reg        [7:0]    io_input_14_delay_15;
  reg        [7:0]    io_input_15_delay_1;
  reg        [7:0]    io_input_15_delay_2;
  reg        [7:0]    io_input_15_delay_3;
  reg        [7:0]    io_input_15_delay_4;
  reg        [7:0]    io_input_15_delay_5;
  reg        [7:0]    io_input_15_delay_6;
  reg        [7:0]    io_input_15_delay_7;
  reg        [7:0]    io_input_15_delay_8;
  reg        [7:0]    io_input_15_delay_9;
  reg        [7:0]    io_input_15_delay_10;
  reg        [7:0]    io_input_15_delay_11;
  reg        [7:0]    io_input_15_delay_12;
  reg        [7:0]    io_input_15_delay_13;
  reg        [7:0]    io_input_15_delay_14;
  reg        [7:0]    io_input_15_delay_15;
  reg        [7:0]    io_input_15_delay_16;

  assign io_output_0 = io_input_0_delay_1;
  assign io_output_1 = io_input_1_delay_2;
  assign io_output_2 = io_input_2_delay_3;
  assign io_output_3 = io_input_3_delay_4;
  assign io_output_4 = io_input_4_delay_5;
  assign io_output_5 = io_input_5_delay_6;
  assign io_output_6 = io_input_6_delay_7;
  assign io_output_7 = io_input_7_delay_8;
  assign io_output_8 = io_input_8_delay_9;
  assign io_output_9 = io_input_9_delay_10;
  assign io_output_10 = io_input_10_delay_11;
  assign io_output_11 = io_input_11_delay_12;
  assign io_output_12 = io_input_12_delay_13;
  assign io_output_13 = io_input_13_delay_14;
  assign io_output_14 = io_input_14_delay_15;
  assign io_output_15 = io_input_15_delay_16;
  always @(posedge clk) begin
    io_input_0_delay_1 <= io_input_0;
    io_input_1_delay_1 <= io_input_1;
    io_input_1_delay_2 <= io_input_1_delay_1;
    io_input_2_delay_1 <= io_input_2;
    io_input_2_delay_2 <= io_input_2_delay_1;
    io_input_2_delay_3 <= io_input_2_delay_2;
    io_input_3_delay_1 <= io_input_3;
    io_input_3_delay_2 <= io_input_3_delay_1;
    io_input_3_delay_3 <= io_input_3_delay_2;
    io_input_3_delay_4 <= io_input_3_delay_3;
    io_input_4_delay_1 <= io_input_4;
    io_input_4_delay_2 <= io_input_4_delay_1;
    io_input_4_delay_3 <= io_input_4_delay_2;
    io_input_4_delay_4 <= io_input_4_delay_3;
    io_input_4_delay_5 <= io_input_4_delay_4;
    io_input_5_delay_1 <= io_input_5;
    io_input_5_delay_2 <= io_input_5_delay_1;
    io_input_5_delay_3 <= io_input_5_delay_2;
    io_input_5_delay_4 <= io_input_5_delay_3;
    io_input_5_delay_5 <= io_input_5_delay_4;
    io_input_5_delay_6 <= io_input_5_delay_5;
    io_input_6_delay_1 <= io_input_6;
    io_input_6_delay_2 <= io_input_6_delay_1;
    io_input_6_delay_3 <= io_input_6_delay_2;
    io_input_6_delay_4 <= io_input_6_delay_3;
    io_input_6_delay_5 <= io_input_6_delay_4;
    io_input_6_delay_6 <= io_input_6_delay_5;
    io_input_6_delay_7 <= io_input_6_delay_6;
    io_input_7_delay_1 <= io_input_7;
    io_input_7_delay_2 <= io_input_7_delay_1;
    io_input_7_delay_3 <= io_input_7_delay_2;
    io_input_7_delay_4 <= io_input_7_delay_3;
    io_input_7_delay_5 <= io_input_7_delay_4;
    io_input_7_delay_6 <= io_input_7_delay_5;
    io_input_7_delay_7 <= io_input_7_delay_6;
    io_input_7_delay_8 <= io_input_7_delay_7;
    io_input_8_delay_1 <= io_input_8;
    io_input_8_delay_2 <= io_input_8_delay_1;
    io_input_8_delay_3 <= io_input_8_delay_2;
    io_input_8_delay_4 <= io_input_8_delay_3;
    io_input_8_delay_5 <= io_input_8_delay_4;
    io_input_8_delay_6 <= io_input_8_delay_5;
    io_input_8_delay_7 <= io_input_8_delay_6;
    io_input_8_delay_8 <= io_input_8_delay_7;
    io_input_8_delay_9 <= io_input_8_delay_8;
    io_input_9_delay_1 <= io_input_9;
    io_input_9_delay_2 <= io_input_9_delay_1;
    io_input_9_delay_3 <= io_input_9_delay_2;
    io_input_9_delay_4 <= io_input_9_delay_3;
    io_input_9_delay_5 <= io_input_9_delay_4;
    io_input_9_delay_6 <= io_input_9_delay_5;
    io_input_9_delay_7 <= io_input_9_delay_6;
    io_input_9_delay_8 <= io_input_9_delay_7;
    io_input_9_delay_9 <= io_input_9_delay_8;
    io_input_9_delay_10 <= io_input_9_delay_9;
    io_input_10_delay_1 <= io_input_10;
    io_input_10_delay_2 <= io_input_10_delay_1;
    io_input_10_delay_3 <= io_input_10_delay_2;
    io_input_10_delay_4 <= io_input_10_delay_3;
    io_input_10_delay_5 <= io_input_10_delay_4;
    io_input_10_delay_6 <= io_input_10_delay_5;
    io_input_10_delay_7 <= io_input_10_delay_6;
    io_input_10_delay_8 <= io_input_10_delay_7;
    io_input_10_delay_9 <= io_input_10_delay_8;
    io_input_10_delay_10 <= io_input_10_delay_9;
    io_input_10_delay_11 <= io_input_10_delay_10;
    io_input_11_delay_1 <= io_input_11;
    io_input_11_delay_2 <= io_input_11_delay_1;
    io_input_11_delay_3 <= io_input_11_delay_2;
    io_input_11_delay_4 <= io_input_11_delay_3;
    io_input_11_delay_5 <= io_input_11_delay_4;
    io_input_11_delay_6 <= io_input_11_delay_5;
    io_input_11_delay_7 <= io_input_11_delay_6;
    io_input_11_delay_8 <= io_input_11_delay_7;
    io_input_11_delay_9 <= io_input_11_delay_8;
    io_input_11_delay_10 <= io_input_11_delay_9;
    io_input_11_delay_11 <= io_input_11_delay_10;
    io_input_11_delay_12 <= io_input_11_delay_11;
    io_input_12_delay_1 <= io_input_12;
    io_input_12_delay_2 <= io_input_12_delay_1;
    io_input_12_delay_3 <= io_input_12_delay_2;
    io_input_12_delay_4 <= io_input_12_delay_3;
    io_input_12_delay_5 <= io_input_12_delay_4;
    io_input_12_delay_6 <= io_input_12_delay_5;
    io_input_12_delay_7 <= io_input_12_delay_6;
    io_input_12_delay_8 <= io_input_12_delay_7;
    io_input_12_delay_9 <= io_input_12_delay_8;
    io_input_12_delay_10 <= io_input_12_delay_9;
    io_input_12_delay_11 <= io_input_12_delay_10;
    io_input_12_delay_12 <= io_input_12_delay_11;
    io_input_12_delay_13 <= io_input_12_delay_12;
    io_input_13_delay_1 <= io_input_13;
    io_input_13_delay_2 <= io_input_13_delay_1;
    io_input_13_delay_3 <= io_input_13_delay_2;
    io_input_13_delay_4 <= io_input_13_delay_3;
    io_input_13_delay_5 <= io_input_13_delay_4;
    io_input_13_delay_6 <= io_input_13_delay_5;
    io_input_13_delay_7 <= io_input_13_delay_6;
    io_input_13_delay_8 <= io_input_13_delay_7;
    io_input_13_delay_9 <= io_input_13_delay_8;
    io_input_13_delay_10 <= io_input_13_delay_9;
    io_input_13_delay_11 <= io_input_13_delay_10;
    io_input_13_delay_12 <= io_input_13_delay_11;
    io_input_13_delay_13 <= io_input_13_delay_12;
    io_input_13_delay_14 <= io_input_13_delay_13;
    io_input_14_delay_1 <= io_input_14;
    io_input_14_delay_2 <= io_input_14_delay_1;
    io_input_14_delay_3 <= io_input_14_delay_2;
    io_input_14_delay_4 <= io_input_14_delay_3;
    io_input_14_delay_5 <= io_input_14_delay_4;
    io_input_14_delay_6 <= io_input_14_delay_5;
    io_input_14_delay_7 <= io_input_14_delay_6;
    io_input_14_delay_8 <= io_input_14_delay_7;
    io_input_14_delay_9 <= io_input_14_delay_8;
    io_input_14_delay_10 <= io_input_14_delay_9;
    io_input_14_delay_11 <= io_input_14_delay_10;
    io_input_14_delay_12 <= io_input_14_delay_11;
    io_input_14_delay_13 <= io_input_14_delay_12;
    io_input_14_delay_14 <= io_input_14_delay_13;
    io_input_14_delay_15 <= io_input_14_delay_14;
    io_input_15_delay_1 <= io_input_15;
    io_input_15_delay_2 <= io_input_15_delay_1;
    io_input_15_delay_3 <= io_input_15_delay_2;
    io_input_15_delay_4 <= io_input_15_delay_3;
    io_input_15_delay_5 <= io_input_15_delay_4;
    io_input_15_delay_6 <= io_input_15_delay_5;
    io_input_15_delay_7 <= io_input_15_delay_6;
    io_input_15_delay_8 <= io_input_15_delay_7;
    io_input_15_delay_9 <= io_input_15_delay_8;
    io_input_15_delay_10 <= io_input_15_delay_9;
    io_input_15_delay_11 <= io_input_15_delay_10;
    io_input_15_delay_12 <= io_input_15_delay_11;
    io_input_15_delay_13 <= io_input_15_delay_12;
    io_input_15_delay_14 <= io_input_15_delay_13;
    io_input_15_delay_15 <= io_input_15_delay_14;
    io_input_15_delay_16 <= io_input_15_delay_15;
  end


endmodule

module ProcessingElement_255 (
  input  wire [7:0]    io_inputA,
  input  wire [7:0]    io_inputB,
  input  wire [19:0]   io_inputC,
  input  wire          io_inputCaptureEnableB,
  output wire [19:0]   io_outputC,
  input  wire          clk,
  input  wire          reset
);

  wire       [19:0]   _zz__zz_io_outputC;
  wire       [15:0]   _zz__zz_io_outputC_1;
  reg        [7:0]    io_inputB_regNextWhen;
  reg        [19:0]   _zz_io_outputC;

  assign _zz__zz_io_outputC_1 = ($signed(io_inputA) * $signed(io_inputB_regNextWhen));
  assign _zz__zz_io_outputC = {{4{_zz__zz_io_outputC_1[15]}}, _zz__zz_io_outputC_1};
  assign io_outputC = _zz_io_outputC;
  always @(posedge clk) begin
    if(reset) begin
      io_inputB_regNextWhen <= 8'h0;
      _zz_io_outputC <= 20'h0;
    end else begin
      if(io_inputCaptureEnableB) begin
        io_inputB_regNextWhen <= io_inputB;
      end
      _zz_io_outputC <= ($signed(_zz__zz_io_outputC) + $signed(io_inputC));
    end
  end


endmodule

//ProcessingElement_254 replaced by ProcessingElement_240

//ProcessingElement_253 replaced by ProcessingElement_240

//ProcessingElement_252 replaced by ProcessingElement_240

//ProcessingElement_251 replaced by ProcessingElement_240

//ProcessingElement_250 replaced by ProcessingElement_240

//ProcessingElement_249 replaced by ProcessingElement_240

//ProcessingElement_248 replaced by ProcessingElement_240

//ProcessingElement_247 replaced by ProcessingElement_240

//ProcessingElement_246 replaced by ProcessingElement_240

//ProcessingElement_245 replaced by ProcessingElement_240

//ProcessingElement_244 replaced by ProcessingElement_240

//ProcessingElement_243 replaced by ProcessingElement_240

//ProcessingElement_242 replaced by ProcessingElement_240

//ProcessingElement_241 replaced by ProcessingElement_240

module ProcessingElement_240 (
  input  wire [7:0]    io_inputA,
  input  wire [7:0]    io_inputB,
  input  wire [19:0]   io_inputC,
  input  wire          io_inputCaptureEnableB,
  output wire [7:0]    io_outputA,
  output wire [19:0]   io_outputC,
  input  wire          clk,
  input  wire          reset
);

  wire       [19:0]   _zz__zz_io_outputC;
  wire       [15:0]   _zz__zz_io_outputC_1;
  reg        [7:0]    io_inputB_regNextWhen;
  reg        [7:0]    io_inputA_regNext;
  reg        [19:0]   _zz_io_outputC;

  assign _zz__zz_io_outputC_1 = ($signed(io_inputA) * $signed(io_inputB_regNextWhen));
  assign _zz__zz_io_outputC = {{4{_zz__zz_io_outputC_1[15]}}, _zz__zz_io_outputC_1};
  assign io_outputA = io_inputA_regNext;
  assign io_outputC = _zz_io_outputC;
  always @(posedge clk) begin
    if(reset) begin
      io_inputB_regNextWhen <= 8'h0;
      io_inputA_regNext <= 8'h0;
      _zz_io_outputC <= 20'h0;
    end else begin
      if(io_inputCaptureEnableB) begin
        io_inputB_regNextWhen <= io_inputB;
      end
      io_inputA_regNext <= io_inputA;
      _zz_io_outputC <= ($signed(_zz__zz_io_outputC) + $signed(io_inputC));
    end
  end


endmodule

//ProcessingElement_239 replaced by ProcessingElement_159

//ProcessingElement_238 replaced by ProcessingElement_144

//ProcessingElement_237 replaced by ProcessingElement_144

//ProcessingElement_236 replaced by ProcessingElement_144

//ProcessingElement_235 replaced by ProcessingElement_144

//ProcessingElement_234 replaced by ProcessingElement_144

//ProcessingElement_233 replaced by ProcessingElement_144

//ProcessingElement_232 replaced by ProcessingElement_144

//ProcessingElement_231 replaced by ProcessingElement_144

//ProcessingElement_230 replaced by ProcessingElement_144

//ProcessingElement_229 replaced by ProcessingElement_144

//ProcessingElement_228 replaced by ProcessingElement_144

//ProcessingElement_227 replaced by ProcessingElement_144

//ProcessingElement_226 replaced by ProcessingElement_144

//ProcessingElement_225 replaced by ProcessingElement_144

//ProcessingElement_224 replaced by ProcessingElement_144

//ProcessingElement_223 replaced by ProcessingElement_159

//ProcessingElement_222 replaced by ProcessingElement_144

//ProcessingElement_221 replaced by ProcessingElement_144

//ProcessingElement_220 replaced by ProcessingElement_144

//ProcessingElement_219 replaced by ProcessingElement_144

//ProcessingElement_218 replaced by ProcessingElement_144

//ProcessingElement_217 replaced by ProcessingElement_144

//ProcessingElement_216 replaced by ProcessingElement_144

//ProcessingElement_215 replaced by ProcessingElement_144

//ProcessingElement_214 replaced by ProcessingElement_144

//ProcessingElement_213 replaced by ProcessingElement_144

//ProcessingElement_212 replaced by ProcessingElement_144

//ProcessingElement_211 replaced by ProcessingElement_144

//ProcessingElement_210 replaced by ProcessingElement_144

//ProcessingElement_209 replaced by ProcessingElement_144

//ProcessingElement_208 replaced by ProcessingElement_144

//ProcessingElement_207 replaced by ProcessingElement_159

//ProcessingElement_206 replaced by ProcessingElement_144

//ProcessingElement_205 replaced by ProcessingElement_144

//ProcessingElement_204 replaced by ProcessingElement_144

//ProcessingElement_203 replaced by ProcessingElement_144

//ProcessingElement_202 replaced by ProcessingElement_144

//ProcessingElement_201 replaced by ProcessingElement_144

//ProcessingElement_200 replaced by ProcessingElement_144

//ProcessingElement_199 replaced by ProcessingElement_144

//ProcessingElement_198 replaced by ProcessingElement_144

//ProcessingElement_197 replaced by ProcessingElement_144

//ProcessingElement_196 replaced by ProcessingElement_144

//ProcessingElement_195 replaced by ProcessingElement_144

//ProcessingElement_194 replaced by ProcessingElement_144

//ProcessingElement_193 replaced by ProcessingElement_144

//ProcessingElement_192 replaced by ProcessingElement_144

//ProcessingElement_191 replaced by ProcessingElement_159

//ProcessingElement_190 replaced by ProcessingElement_144

//ProcessingElement_189 replaced by ProcessingElement_144

//ProcessingElement_188 replaced by ProcessingElement_144

//ProcessingElement_187 replaced by ProcessingElement_144

//ProcessingElement_186 replaced by ProcessingElement_144

//ProcessingElement_185 replaced by ProcessingElement_144

//ProcessingElement_184 replaced by ProcessingElement_144

//ProcessingElement_183 replaced by ProcessingElement_144

//ProcessingElement_182 replaced by ProcessingElement_144

//ProcessingElement_181 replaced by ProcessingElement_144

//ProcessingElement_180 replaced by ProcessingElement_144

//ProcessingElement_179 replaced by ProcessingElement_144

//ProcessingElement_178 replaced by ProcessingElement_144

//ProcessingElement_177 replaced by ProcessingElement_144

//ProcessingElement_176 replaced by ProcessingElement_144

//ProcessingElement_175 replaced by ProcessingElement_159

//ProcessingElement_174 replaced by ProcessingElement_144

//ProcessingElement_173 replaced by ProcessingElement_144

//ProcessingElement_172 replaced by ProcessingElement_144

//ProcessingElement_171 replaced by ProcessingElement_144

//ProcessingElement_170 replaced by ProcessingElement_144

//ProcessingElement_169 replaced by ProcessingElement_144

//ProcessingElement_168 replaced by ProcessingElement_144

//ProcessingElement_167 replaced by ProcessingElement_144

//ProcessingElement_166 replaced by ProcessingElement_144

//ProcessingElement_165 replaced by ProcessingElement_144

//ProcessingElement_164 replaced by ProcessingElement_144

//ProcessingElement_163 replaced by ProcessingElement_144

//ProcessingElement_162 replaced by ProcessingElement_144

//ProcessingElement_161 replaced by ProcessingElement_144

//ProcessingElement_160 replaced by ProcessingElement_144

module ProcessingElement_159 (
  input  wire [7:0]    io_inputA,
  input  wire [7:0]    io_inputB,
  input  wire [19:0]   io_inputC,
  input  wire          io_inputCaptureEnableB,
  output wire [7:0]    io_outputB,
  output wire [19:0]   io_outputC,
  input  wire          clk,
  input  wire          reset
);

  wire       [19:0]   _zz__zz_io_outputC;
  wire       [15:0]   _zz__zz_io_outputC_1;
  reg        [7:0]    io_inputB_regNextWhen;
  reg        [19:0]   _zz_io_outputC;

  assign _zz__zz_io_outputC_1 = ($signed(io_inputA) * $signed(io_inputB_regNextWhen));
  assign _zz__zz_io_outputC = {{4{_zz__zz_io_outputC_1[15]}}, _zz__zz_io_outputC_1};
  assign io_outputB = io_inputB_regNextWhen;
  assign io_outputC = _zz_io_outputC;
  always @(posedge clk) begin
    if(reset) begin
      io_inputB_regNextWhen <= 8'h0;
      _zz_io_outputC <= 20'h0;
    end else begin
      if(io_inputCaptureEnableB) begin
        io_inputB_regNextWhen <= io_inputB;
      end
      _zz_io_outputC <= ($signed(_zz__zz_io_outputC) + $signed(io_inputC));
    end
  end


endmodule

//ProcessingElement_158 replaced by ProcessingElement_144

//ProcessingElement_157 replaced by ProcessingElement_144

//ProcessingElement_156 replaced by ProcessingElement_144

//ProcessingElement_155 replaced by ProcessingElement_144

//ProcessingElement_154 replaced by ProcessingElement_144

//ProcessingElement_153 replaced by ProcessingElement_144

//ProcessingElement_152 replaced by ProcessingElement_144

//ProcessingElement_151 replaced by ProcessingElement_144

//ProcessingElement_150 replaced by ProcessingElement_144

//ProcessingElement_149 replaced by ProcessingElement_144

//ProcessingElement_148 replaced by ProcessingElement_144

//ProcessingElement_147 replaced by ProcessingElement_144

//ProcessingElement_146 replaced by ProcessingElement_144

//ProcessingElement_145 replaced by ProcessingElement_144

module ProcessingElement_144 (
  input  wire [7:0]    io_inputA,
  input  wire [7:0]    io_inputB,
  input  wire [19:0]   io_inputC,
  input  wire          io_inputCaptureEnableB,
  output wire [7:0]    io_outputA,
  output wire [7:0]    io_outputB,
  output wire [19:0]   io_outputC,
  input  wire          clk,
  input  wire          reset
);

  wire       [19:0]   _zz__zz_io_outputC;
  wire       [15:0]   _zz__zz_io_outputC_1;
  reg        [7:0]    io_inputB_regNextWhen;
  reg        [7:0]    io_inputA_regNext;
  reg        [19:0]   _zz_io_outputC;

  assign _zz__zz_io_outputC_1 = ($signed(io_inputA) * $signed(io_inputB_regNextWhen));
  assign _zz__zz_io_outputC = {{4{_zz__zz_io_outputC_1[15]}}, _zz__zz_io_outputC_1};
  assign io_outputA = io_inputA_regNext;
  assign io_outputB = io_inputB_regNextWhen;
  assign io_outputC = _zz_io_outputC;
  always @(posedge clk) begin
    if(reset) begin
      io_inputB_regNextWhen <= 8'h0;
      io_inputA_regNext <= 8'h0;
      _zz_io_outputC <= 20'h0;
    end else begin
      if(io_inputCaptureEnableB) begin
        io_inputB_regNextWhen <= io_inputB;
      end
      io_inputA_regNext <= io_inputA;
      _zz_io_outputC <= ($signed(_zz__zz_io_outputC) + $signed(io_inputC));
    end
  end


endmodule

module ProcessingElement_143 (
  input  wire [7:0]    io_inputA,
  input  wire [7:0]    io_inputB,
  input  wire [18:0]   io_inputC,
  input  wire          io_inputCaptureEnableB,
  output wire [7:0]    io_outputB,
  output wire [19:0]   io_outputC,
  input  wire          clk,
  input  wire          reset
);

  wire       [18:0]   _zz__zz_io_outputC;
  wire       [18:0]   _zz__zz_io_outputC_1;
  wire       [15:0]   _zz__zz_io_outputC_2;
  reg        [7:0]    io_inputB_regNextWhen;
  reg        [19:0]   _zz_io_outputC;

  assign _zz__zz_io_outputC = ($signed(_zz__zz_io_outputC_1) + $signed(io_inputC));
  assign _zz__zz_io_outputC_2 = ($signed(io_inputA) * $signed(io_inputB_regNextWhen));
  assign _zz__zz_io_outputC_1 = {{3{_zz__zz_io_outputC_2[15]}}, _zz__zz_io_outputC_2};
  assign io_outputB = io_inputB_regNextWhen;
  assign io_outputC = _zz_io_outputC;
  always @(posedge clk) begin
    if(reset) begin
      io_inputB_regNextWhen <= 8'h0;
      _zz_io_outputC <= 20'h0;
    end else begin
      if(io_inputCaptureEnableB) begin
        io_inputB_regNextWhen <= io_inputB;
      end
      _zz_io_outputC <= {{1{_zz__zz_io_outputC[18]}}, _zz__zz_io_outputC};
    end
  end


endmodule

//ProcessingElement_142 replaced by ProcessingElement_128

//ProcessingElement_141 replaced by ProcessingElement_128

//ProcessingElement_140 replaced by ProcessingElement_128

//ProcessingElement_139 replaced by ProcessingElement_128

//ProcessingElement_138 replaced by ProcessingElement_128

//ProcessingElement_137 replaced by ProcessingElement_128

//ProcessingElement_136 replaced by ProcessingElement_128

//ProcessingElement_135 replaced by ProcessingElement_128

//ProcessingElement_134 replaced by ProcessingElement_128

//ProcessingElement_133 replaced by ProcessingElement_128

//ProcessingElement_132 replaced by ProcessingElement_128

//ProcessingElement_131 replaced by ProcessingElement_128

//ProcessingElement_130 replaced by ProcessingElement_128

//ProcessingElement_129 replaced by ProcessingElement_128

module ProcessingElement_128 (
  input  wire [7:0]    io_inputA,
  input  wire [7:0]    io_inputB,
  input  wire [18:0]   io_inputC,
  input  wire          io_inputCaptureEnableB,
  output wire [7:0]    io_outputA,
  output wire [7:0]    io_outputB,
  output wire [19:0]   io_outputC,
  input  wire          clk,
  input  wire          reset
);

  wire       [18:0]   _zz__zz_io_outputC;
  wire       [18:0]   _zz__zz_io_outputC_1;
  wire       [15:0]   _zz__zz_io_outputC_2;
  reg        [7:0]    io_inputB_regNextWhen;
  reg        [7:0]    io_inputA_regNext;
  reg        [19:0]   _zz_io_outputC;

  assign _zz__zz_io_outputC = ($signed(_zz__zz_io_outputC_1) + $signed(io_inputC));
  assign _zz__zz_io_outputC_2 = ($signed(io_inputA) * $signed(io_inputB_regNextWhen));
  assign _zz__zz_io_outputC_1 = {{3{_zz__zz_io_outputC_2[15]}}, _zz__zz_io_outputC_2};
  assign io_outputA = io_inputA_regNext;
  assign io_outputB = io_inputB_regNextWhen;
  assign io_outputC = _zz_io_outputC;
  always @(posedge clk) begin
    if(reset) begin
      io_inputB_regNextWhen <= 8'h0;
      io_inputA_regNext <= 8'h0;
      _zz_io_outputC <= 20'h0;
    end else begin
      if(io_inputCaptureEnableB) begin
        io_inputB_regNextWhen <= io_inputB;
      end
      io_inputA_regNext <= io_inputA;
      _zz_io_outputC <= {{1{_zz__zz_io_outputC[18]}}, _zz__zz_io_outputC};
    end
  end


endmodule

//ProcessingElement_127 replaced by ProcessingElement_95

//ProcessingElement_126 replaced by ProcessingElement_80

//ProcessingElement_125 replaced by ProcessingElement_80

//ProcessingElement_124 replaced by ProcessingElement_80

//ProcessingElement_123 replaced by ProcessingElement_80

//ProcessingElement_122 replaced by ProcessingElement_80

//ProcessingElement_121 replaced by ProcessingElement_80

//ProcessingElement_120 replaced by ProcessingElement_80

//ProcessingElement_119 replaced by ProcessingElement_80

//ProcessingElement_118 replaced by ProcessingElement_80

//ProcessingElement_117 replaced by ProcessingElement_80

//ProcessingElement_116 replaced by ProcessingElement_80

//ProcessingElement_115 replaced by ProcessingElement_80

//ProcessingElement_114 replaced by ProcessingElement_80

//ProcessingElement_113 replaced by ProcessingElement_80

//ProcessingElement_112 replaced by ProcessingElement_80

//ProcessingElement_111 replaced by ProcessingElement_95

//ProcessingElement_110 replaced by ProcessingElement_80

//ProcessingElement_109 replaced by ProcessingElement_80

//ProcessingElement_108 replaced by ProcessingElement_80

//ProcessingElement_107 replaced by ProcessingElement_80

//ProcessingElement_106 replaced by ProcessingElement_80

//ProcessingElement_105 replaced by ProcessingElement_80

//ProcessingElement_104 replaced by ProcessingElement_80

//ProcessingElement_103 replaced by ProcessingElement_80

//ProcessingElement_102 replaced by ProcessingElement_80

//ProcessingElement_101 replaced by ProcessingElement_80

//ProcessingElement_100 replaced by ProcessingElement_80

//ProcessingElement_99 replaced by ProcessingElement_80

//ProcessingElement_98 replaced by ProcessingElement_80

//ProcessingElement_97 replaced by ProcessingElement_80

//ProcessingElement_96 replaced by ProcessingElement_80

module ProcessingElement_95 (
  input  wire [7:0]    io_inputA,
  input  wire [7:0]    io_inputB,
  input  wire [18:0]   io_inputC,
  input  wire          io_inputCaptureEnableB,
  output wire [7:0]    io_outputB,
  output wire [18:0]   io_outputC,
  input  wire          clk,
  input  wire          reset
);

  wire       [18:0]   _zz__zz_io_outputC;
  wire       [15:0]   _zz__zz_io_outputC_1;
  reg        [7:0]    io_inputB_regNextWhen;
  reg        [18:0]   _zz_io_outputC;

  assign _zz__zz_io_outputC_1 = ($signed(io_inputA) * $signed(io_inputB_regNextWhen));
  assign _zz__zz_io_outputC = {{3{_zz__zz_io_outputC_1[15]}}, _zz__zz_io_outputC_1};
  assign io_outputB = io_inputB_regNextWhen;
  assign io_outputC = _zz_io_outputC;
  always @(posedge clk) begin
    if(reset) begin
      io_inputB_regNextWhen <= 8'h0;
      _zz_io_outputC <= 19'h0;
    end else begin
      if(io_inputCaptureEnableB) begin
        io_inputB_regNextWhen <= io_inputB;
      end
      _zz_io_outputC <= ($signed(_zz__zz_io_outputC) + $signed(io_inputC));
    end
  end


endmodule

//ProcessingElement_94 replaced by ProcessingElement_80

//ProcessingElement_93 replaced by ProcessingElement_80

//ProcessingElement_92 replaced by ProcessingElement_80

//ProcessingElement_91 replaced by ProcessingElement_80

//ProcessingElement_90 replaced by ProcessingElement_80

//ProcessingElement_89 replaced by ProcessingElement_80

//ProcessingElement_88 replaced by ProcessingElement_80

//ProcessingElement_87 replaced by ProcessingElement_80

//ProcessingElement_86 replaced by ProcessingElement_80

//ProcessingElement_85 replaced by ProcessingElement_80

//ProcessingElement_84 replaced by ProcessingElement_80

//ProcessingElement_83 replaced by ProcessingElement_80

//ProcessingElement_82 replaced by ProcessingElement_80

//ProcessingElement_81 replaced by ProcessingElement_80

module ProcessingElement_80 (
  input  wire [7:0]    io_inputA,
  input  wire [7:0]    io_inputB,
  input  wire [18:0]   io_inputC,
  input  wire          io_inputCaptureEnableB,
  output wire [7:0]    io_outputA,
  output wire [7:0]    io_outputB,
  output wire [18:0]   io_outputC,
  input  wire          clk,
  input  wire          reset
);

  wire       [18:0]   _zz__zz_io_outputC;
  wire       [15:0]   _zz__zz_io_outputC_1;
  reg        [7:0]    io_inputB_regNextWhen;
  reg        [7:0]    io_inputA_regNext;
  reg        [18:0]   _zz_io_outputC;

  assign _zz__zz_io_outputC_1 = ($signed(io_inputA) * $signed(io_inputB_regNextWhen));
  assign _zz__zz_io_outputC = {{3{_zz__zz_io_outputC_1[15]}}, _zz__zz_io_outputC_1};
  assign io_outputA = io_inputA_regNext;
  assign io_outputB = io_inputB_regNextWhen;
  assign io_outputC = _zz_io_outputC;
  always @(posedge clk) begin
    if(reset) begin
      io_inputB_regNextWhen <= 8'h0;
      io_inputA_regNext <= 8'h0;
      _zz_io_outputC <= 19'h0;
    end else begin
      if(io_inputCaptureEnableB) begin
        io_inputB_regNextWhen <= io_inputB;
      end
      io_inputA_regNext <= io_inputA;
      _zz_io_outputC <= ($signed(_zz__zz_io_outputC) + $signed(io_inputC));
    end
  end


endmodule

module ProcessingElement_79 (
  input  wire [7:0]    io_inputA,
  input  wire [7:0]    io_inputB,
  input  wire [17:0]   io_inputC,
  input  wire          io_inputCaptureEnableB,
  output wire [7:0]    io_outputB,
  output wire [18:0]   io_outputC,
  input  wire          clk,
  input  wire          reset
);

  wire       [17:0]   _zz__zz_io_outputC;
  wire       [17:0]   _zz__zz_io_outputC_1;
  wire       [15:0]   _zz__zz_io_outputC_2;
  reg        [7:0]    io_inputB_regNextWhen;
  reg        [18:0]   _zz_io_outputC;

  assign _zz__zz_io_outputC = ($signed(_zz__zz_io_outputC_1) + $signed(io_inputC));
  assign _zz__zz_io_outputC_2 = ($signed(io_inputA) * $signed(io_inputB_regNextWhen));
  assign _zz__zz_io_outputC_1 = {{2{_zz__zz_io_outputC_2[15]}}, _zz__zz_io_outputC_2};
  assign io_outputB = io_inputB_regNextWhen;
  assign io_outputC = _zz_io_outputC;
  always @(posedge clk) begin
    if(reset) begin
      io_inputB_regNextWhen <= 8'h0;
      _zz_io_outputC <= 19'h0;
    end else begin
      if(io_inputCaptureEnableB) begin
        io_inputB_regNextWhen <= io_inputB;
      end
      _zz_io_outputC <= {{1{_zz__zz_io_outputC[17]}}, _zz__zz_io_outputC};
    end
  end


endmodule

//ProcessingElement_78 replaced by ProcessingElement_64

//ProcessingElement_77 replaced by ProcessingElement_64

//ProcessingElement_76 replaced by ProcessingElement_64

//ProcessingElement_75 replaced by ProcessingElement_64

//ProcessingElement_74 replaced by ProcessingElement_64

//ProcessingElement_73 replaced by ProcessingElement_64

//ProcessingElement_72 replaced by ProcessingElement_64

//ProcessingElement_71 replaced by ProcessingElement_64

//ProcessingElement_70 replaced by ProcessingElement_64

//ProcessingElement_69 replaced by ProcessingElement_64

//ProcessingElement_68 replaced by ProcessingElement_64

//ProcessingElement_67 replaced by ProcessingElement_64

//ProcessingElement_66 replaced by ProcessingElement_64

//ProcessingElement_65 replaced by ProcessingElement_64

module ProcessingElement_64 (
  input  wire [7:0]    io_inputA,
  input  wire [7:0]    io_inputB,
  input  wire [17:0]   io_inputC,
  input  wire          io_inputCaptureEnableB,
  output wire [7:0]    io_outputA,
  output wire [7:0]    io_outputB,
  output wire [18:0]   io_outputC,
  input  wire          clk,
  input  wire          reset
);

  wire       [17:0]   _zz__zz_io_outputC;
  wire       [17:0]   _zz__zz_io_outputC_1;
  wire       [15:0]   _zz__zz_io_outputC_2;
  reg        [7:0]    io_inputB_regNextWhen;
  reg        [7:0]    io_inputA_regNext;
  reg        [18:0]   _zz_io_outputC;

  assign _zz__zz_io_outputC = ($signed(_zz__zz_io_outputC_1) + $signed(io_inputC));
  assign _zz__zz_io_outputC_2 = ($signed(io_inputA) * $signed(io_inputB_regNextWhen));
  assign _zz__zz_io_outputC_1 = {{2{_zz__zz_io_outputC_2[15]}}, _zz__zz_io_outputC_2};
  assign io_outputA = io_inputA_regNext;
  assign io_outputB = io_inputB_regNextWhen;
  assign io_outputC = _zz_io_outputC;
  always @(posedge clk) begin
    if(reset) begin
      io_inputB_regNextWhen <= 8'h0;
      io_inputA_regNext <= 8'h0;
      _zz_io_outputC <= 19'h0;
    end else begin
      if(io_inputCaptureEnableB) begin
        io_inputB_regNextWhen <= io_inputB;
      end
      io_inputA_regNext <= io_inputA;
      _zz_io_outputC <= {{1{_zz__zz_io_outputC[17]}}, _zz__zz_io_outputC};
    end
  end


endmodule

module ProcessingElement_63 (
  input  wire [7:0]    io_inputA,
  input  wire [7:0]    io_inputB,
  input  wire [17:0]   io_inputC,
  input  wire          io_inputCaptureEnableB,
  output wire [7:0]    io_outputB,
  output wire [17:0]   io_outputC,
  input  wire          clk,
  input  wire          reset
);

  wire       [17:0]   _zz__zz_io_outputC;
  wire       [15:0]   _zz__zz_io_outputC_1;
  reg        [7:0]    io_inputB_regNextWhen;
  reg        [17:0]   _zz_io_outputC;

  assign _zz__zz_io_outputC_1 = ($signed(io_inputA) * $signed(io_inputB_regNextWhen));
  assign _zz__zz_io_outputC = {{2{_zz__zz_io_outputC_1[15]}}, _zz__zz_io_outputC_1};
  assign io_outputB = io_inputB_regNextWhen;
  assign io_outputC = _zz_io_outputC;
  always @(posedge clk) begin
    if(reset) begin
      io_inputB_regNextWhen <= 8'h0;
      _zz_io_outputC <= 18'h0;
    end else begin
      if(io_inputCaptureEnableB) begin
        io_inputB_regNextWhen <= io_inputB;
      end
      _zz_io_outputC <= ($signed(_zz__zz_io_outputC) + $signed(io_inputC));
    end
  end


endmodule

//ProcessingElement_62 replaced by ProcessingElement_48

//ProcessingElement_61 replaced by ProcessingElement_48

//ProcessingElement_60 replaced by ProcessingElement_48

//ProcessingElement_59 replaced by ProcessingElement_48

//ProcessingElement_58 replaced by ProcessingElement_48

//ProcessingElement_57 replaced by ProcessingElement_48

//ProcessingElement_56 replaced by ProcessingElement_48

//ProcessingElement_55 replaced by ProcessingElement_48

//ProcessingElement_54 replaced by ProcessingElement_48

//ProcessingElement_53 replaced by ProcessingElement_48

//ProcessingElement_52 replaced by ProcessingElement_48

//ProcessingElement_51 replaced by ProcessingElement_48

//ProcessingElement_50 replaced by ProcessingElement_48

//ProcessingElement_49 replaced by ProcessingElement_48

module ProcessingElement_48 (
  input  wire [7:0]    io_inputA,
  input  wire [7:0]    io_inputB,
  input  wire [17:0]   io_inputC,
  input  wire          io_inputCaptureEnableB,
  output wire [7:0]    io_outputA,
  output wire [7:0]    io_outputB,
  output wire [17:0]   io_outputC,
  input  wire          clk,
  input  wire          reset
);

  wire       [17:0]   _zz__zz_io_outputC;
  wire       [15:0]   _zz__zz_io_outputC_1;
  reg        [7:0]    io_inputB_regNextWhen;
  reg        [7:0]    io_inputA_regNext;
  reg        [17:0]   _zz_io_outputC;

  assign _zz__zz_io_outputC_1 = ($signed(io_inputA) * $signed(io_inputB_regNextWhen));
  assign _zz__zz_io_outputC = {{2{_zz__zz_io_outputC_1[15]}}, _zz__zz_io_outputC_1};
  assign io_outputA = io_inputA_regNext;
  assign io_outputB = io_inputB_regNextWhen;
  assign io_outputC = _zz_io_outputC;
  always @(posedge clk) begin
    if(reset) begin
      io_inputB_regNextWhen <= 8'h0;
      io_inputA_regNext <= 8'h0;
      _zz_io_outputC <= 18'h0;
    end else begin
      if(io_inputCaptureEnableB) begin
        io_inputB_regNextWhen <= io_inputB;
      end
      io_inputA_regNext <= io_inputA;
      _zz_io_outputC <= ($signed(_zz__zz_io_outputC) + $signed(io_inputC));
    end
  end


endmodule

module ProcessingElement_47 (
  input  wire [7:0]    io_inputA,
  input  wire [7:0]    io_inputB,
  input  wire [16:0]   io_inputC,
  input  wire          io_inputCaptureEnableB,
  output wire [7:0]    io_outputB,
  output wire [17:0]   io_outputC,
  input  wire          clk,
  input  wire          reset
);

  wire       [16:0]   _zz__zz_io_outputC;
  wire       [16:0]   _zz__zz_io_outputC_1;
  wire       [15:0]   _zz__zz_io_outputC_2;
  reg        [7:0]    io_inputB_regNextWhen;
  reg        [17:0]   _zz_io_outputC;

  assign _zz__zz_io_outputC = ($signed(_zz__zz_io_outputC_1) + $signed(io_inputC));
  assign _zz__zz_io_outputC_2 = ($signed(io_inputA) * $signed(io_inputB_regNextWhen));
  assign _zz__zz_io_outputC_1 = {{1{_zz__zz_io_outputC_2[15]}}, _zz__zz_io_outputC_2};
  assign io_outputB = io_inputB_regNextWhen;
  assign io_outputC = _zz_io_outputC;
  always @(posedge clk) begin
    if(reset) begin
      io_inputB_regNextWhen <= 8'h0;
      _zz_io_outputC <= 18'h0;
    end else begin
      if(io_inputCaptureEnableB) begin
        io_inputB_regNextWhen <= io_inputB;
      end
      _zz_io_outputC <= {{1{_zz__zz_io_outputC[16]}}, _zz__zz_io_outputC};
    end
  end


endmodule

//ProcessingElement_46 replaced by ProcessingElement_32

//ProcessingElement_45 replaced by ProcessingElement_32

//ProcessingElement_44 replaced by ProcessingElement_32

//ProcessingElement_43 replaced by ProcessingElement_32

//ProcessingElement_42 replaced by ProcessingElement_32

//ProcessingElement_41 replaced by ProcessingElement_32

//ProcessingElement_40 replaced by ProcessingElement_32

//ProcessingElement_39 replaced by ProcessingElement_32

//ProcessingElement_38 replaced by ProcessingElement_32

//ProcessingElement_37 replaced by ProcessingElement_32

//ProcessingElement_36 replaced by ProcessingElement_32

//ProcessingElement_35 replaced by ProcessingElement_32

//ProcessingElement_34 replaced by ProcessingElement_32

//ProcessingElement_33 replaced by ProcessingElement_32

module ProcessingElement_32 (
  input  wire [7:0]    io_inputA,
  input  wire [7:0]    io_inputB,
  input  wire [16:0]   io_inputC,
  input  wire          io_inputCaptureEnableB,
  output wire [7:0]    io_outputA,
  output wire [7:0]    io_outputB,
  output wire [17:0]   io_outputC,
  input  wire          clk,
  input  wire          reset
);

  wire       [16:0]   _zz__zz_io_outputC;
  wire       [16:0]   _zz__zz_io_outputC_1;
  wire       [15:0]   _zz__zz_io_outputC_2;
  reg        [7:0]    io_inputB_regNextWhen;
  reg        [7:0]    io_inputA_regNext;
  reg        [17:0]   _zz_io_outputC;

  assign _zz__zz_io_outputC = ($signed(_zz__zz_io_outputC_1) + $signed(io_inputC));
  assign _zz__zz_io_outputC_2 = ($signed(io_inputA) * $signed(io_inputB_regNextWhen));
  assign _zz__zz_io_outputC_1 = {{1{_zz__zz_io_outputC_2[15]}}, _zz__zz_io_outputC_2};
  assign io_outputA = io_inputA_regNext;
  assign io_outputB = io_inputB_regNextWhen;
  assign io_outputC = _zz_io_outputC;
  always @(posedge clk) begin
    if(reset) begin
      io_inputB_regNextWhen <= 8'h0;
      io_inputA_regNext <= 8'h0;
      _zz_io_outputC <= 18'h0;
    end else begin
      if(io_inputCaptureEnableB) begin
        io_inputB_regNextWhen <= io_inputB;
      end
      io_inputA_regNext <= io_inputA;
      _zz_io_outputC <= {{1{_zz__zz_io_outputC[16]}}, _zz__zz_io_outputC};
    end
  end


endmodule

module ProcessingElement_31 (
  input  wire [7:0]    io_inputA,
  input  wire [7:0]    io_inputB,
  input  wire [15:0]   io_inputC,
  input  wire          io_inputCaptureEnableB,
  output wire [7:0]    io_outputB,
  output wire [16:0]   io_outputC,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz_io_outputC;
  wire       [15:0]   _zz__zz_io_outputC_1;
  reg        [7:0]    io_inputB_regNextWhen;
  reg        [16:0]   _zz_io_outputC;

  assign _zz__zz_io_outputC = ($signed(_zz__zz_io_outputC_1) + $signed(io_inputC));
  assign _zz__zz_io_outputC_1 = ($signed(io_inputA) * $signed(io_inputB_regNextWhen));
  assign io_outputB = io_inputB_regNextWhen;
  assign io_outputC = _zz_io_outputC;
  always @(posedge clk) begin
    if(reset) begin
      io_inputB_regNextWhen <= 8'h0;
      _zz_io_outputC <= 17'h0;
    end else begin
      if(io_inputCaptureEnableB) begin
        io_inputB_regNextWhen <= io_inputB;
      end
      _zz_io_outputC <= {{1{_zz__zz_io_outputC[15]}}, _zz__zz_io_outputC};
    end
  end


endmodule

//ProcessingElement_30 replaced by ProcessingElement_16

//ProcessingElement_29 replaced by ProcessingElement_16

//ProcessingElement_28 replaced by ProcessingElement_16

//ProcessingElement_27 replaced by ProcessingElement_16

//ProcessingElement_26 replaced by ProcessingElement_16

//ProcessingElement_25 replaced by ProcessingElement_16

//ProcessingElement_24 replaced by ProcessingElement_16

//ProcessingElement_23 replaced by ProcessingElement_16

//ProcessingElement_22 replaced by ProcessingElement_16

//ProcessingElement_21 replaced by ProcessingElement_16

//ProcessingElement_20 replaced by ProcessingElement_16

//ProcessingElement_19 replaced by ProcessingElement_16

//ProcessingElement_18 replaced by ProcessingElement_16

//ProcessingElement_17 replaced by ProcessingElement_16

module ProcessingElement_16 (
  input  wire [7:0]    io_inputA,
  input  wire [7:0]    io_inputB,
  input  wire [15:0]   io_inputC,
  input  wire          io_inputCaptureEnableB,
  output wire [7:0]    io_outputA,
  output wire [7:0]    io_outputB,
  output wire [16:0]   io_outputC,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz_io_outputC;
  wire       [15:0]   _zz__zz_io_outputC_1;
  reg        [7:0]    io_inputB_regNextWhen;
  reg        [7:0]    io_inputA_regNext;
  reg        [16:0]   _zz_io_outputC;

  assign _zz__zz_io_outputC = ($signed(_zz__zz_io_outputC_1) + $signed(io_inputC));
  assign _zz__zz_io_outputC_1 = ($signed(io_inputA) * $signed(io_inputB_regNextWhen));
  assign io_outputA = io_inputA_regNext;
  assign io_outputB = io_inputB_regNextWhen;
  assign io_outputC = _zz_io_outputC;
  always @(posedge clk) begin
    if(reset) begin
      io_inputB_regNextWhen <= 8'h0;
      io_inputA_regNext <= 8'h0;
      _zz_io_outputC <= 17'h0;
    end else begin
      if(io_inputCaptureEnableB) begin
        io_inputB_regNextWhen <= io_inputB;
      end
      io_inputA_regNext <= io_inputA;
      _zz_io_outputC <= {{1{_zz__zz_io_outputC[15]}}, _zz__zz_io_outputC};
    end
  end


endmodule

module ProcessingElement_15 (
  input  wire [7:0]    io_inputA,
  input  wire [7:0]    io_inputB,
  input  wire          io_inputCaptureEnableB,
  output wire [7:0]    io_outputB,
  output wire [15:0]   io_outputC,
  input  wire          clk,
  input  wire          reset
);

  reg        [7:0]    io_inputB_regNextWhen;
  reg        [15:0]   _zz_io_outputC;

  assign io_outputB = io_inputB_regNextWhen;
  assign io_outputC = _zz_io_outputC;
  always @(posedge clk) begin
    if(reset) begin
      io_inputB_regNextWhen <= 8'h0;
      _zz_io_outputC <= 16'h0;
    end else begin
      if(io_inputCaptureEnableB) begin
        io_inputB_regNextWhen <= io_inputB;
      end
      _zz_io_outputC <= ($signed(io_inputA) * $signed(io_inputB_regNextWhen));
    end
  end


endmodule

//ProcessingElement_14 replaced by ProcessingElement

//ProcessingElement_13 replaced by ProcessingElement

//ProcessingElement_12 replaced by ProcessingElement

//ProcessingElement_11 replaced by ProcessingElement

//ProcessingElement_10 replaced by ProcessingElement

//ProcessingElement_9 replaced by ProcessingElement

//ProcessingElement_8 replaced by ProcessingElement

//ProcessingElement_7 replaced by ProcessingElement

//ProcessingElement_6 replaced by ProcessingElement

//ProcessingElement_5 replaced by ProcessingElement

//ProcessingElement_4 replaced by ProcessingElement

//ProcessingElement_3 replaced by ProcessingElement

//ProcessingElement_2 replaced by ProcessingElement

//ProcessingElement_1 replaced by ProcessingElement

module ProcessingElement (
  input  wire [7:0]    io_inputA,
  input  wire [7:0]    io_inputB,
  input  wire          io_inputCaptureEnableB,
  output wire [7:0]    io_outputA,
  output wire [7:0]    io_outputB,
  output wire [15:0]   io_outputC,
  input  wire          clk,
  input  wire          reset
);

  reg        [7:0]    io_inputB_regNextWhen;
  reg        [7:0]    io_inputA_regNext;
  reg        [15:0]   _zz_io_outputC;

  assign io_outputA = io_inputA_regNext;
  assign io_outputB = io_inputB_regNextWhen;
  assign io_outputC = _zz_io_outputC;
  always @(posedge clk) begin
    if(reset) begin
      io_inputB_regNextWhen <= 8'h0;
      io_inputA_regNext <= 8'h0;
      _zz_io_outputC <= 16'h0;
    end else begin
      if(io_inputCaptureEnableB) begin
        io_inputB_regNextWhen <= io_inputB;
      end
      io_inputA_regNext <= io_inputA;
      _zz_io_outputC <= ($signed(io_inputA) * $signed(io_inputB_regNextWhen));
    end
  end


endmodule
